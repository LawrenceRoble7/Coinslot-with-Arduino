PK   �
.Xƨ�mL  1�     cirkitFile.json�]ێ#7��CƼ)�/��`����>�3���Z�Tn{�������%S*��BeH�R�b��H#����C&��l�~��e����o~�[mֳ7T�gܶ��ο%�٧�z��,ݺOfo������|Qm>~ڬ�z���RS���5���)i��2^U�J�<Y�ٛ_�{�*˦�e;b��5��9��Z�K�B����ƾ.�ڳ�mAjYX�y��/�H�${���<)8��)k�f��D�4�K��bzV�����3����6�`q��)�y��;�E]RQ&��{_��{lQ
mC߈�S"���.jg�p55)ʺ$�t���w-Eh��Y$z�k��F���ʇ��0�7��B����q��2�2�C@��0=��Y'z���*��BR�a�*a��,��*˵����M�g�ʪ6��R��Lfq a�V���t��m�gʈ�.,9�����Ye�Ue����8kS�;A�ʐ�9��@����
�^#ۧ@/�L](]��΂����(K�y�$ �g�K��"�ː�eH�2$t�	]��.("��ўA�G�z�r��e���ZmIM!2�j��BxRǼ�R^�Շ1�SmA�S�����!8�C�T̫JZZ҄�@�y��T]��X�]C�Ι^K�yQS'C�Z���S��ܗ\ٺj(.�M�Pϩl�a����M���^	@���yz ��TbD8�x੮�TM�H"Dϩ�B�sj~ 
�g�D�������gT��Ǘ\c�����b@��R\ 0�B��AD�� H� 4���+0~	���N��!47�/��%L�:mrA������S��fn* 2���N�L�^f@6�5M�M ��y�Tנ�<=;@��s�<�!�u0 �l���S u�˗�~w�y�l��ݳ�������w=�ZT�"B
�R������D<J!$-�כA
�"�d�RZ����tQJ�r�7)r
uН�˨��z�zcQv1QJYW�iRl;FR��bP�	�y�KY1y�5y��<bT1:���:��a��<^/�Y&��,�Y�<(fyP�򠘙�0�Y�A��<�ys>eb�NW)t*:��@]6t7)�����[�,��ty���E�=p�'��əݑɠ��<��d�2��.D)t*ˀ�\�J�g�¦�(wY(��Aʤ]����	J�OxL ϞAʤ]��y)t*����WX(�}Y
���l(�|9сRǗ�.���DP28���(J_f��4o]��=�����{,������{@��x)4��E
��&_�R&�&_�R��Ed�"�HQY��,RL)6�2�7zi��<��y L� ��0̓a��4�Y�L>8�Y�<(fyP���A1˃b��<�y�L��$���+^ʤe��+^J�LNn0�zQ
�|�K����+^J]�s(���2�0�zQ
�|�K�#0����G�I���׋R��+^ʤ]��+^ʴ߅��x)�v��x)����W��I]��+^J]&�&_�R&�L��L�F0���r��}����?�{]���go8��>��~����*_/W��f[����/��iՐ��B�:,��	�W�ec(e��JT�����b^�EE���S1X�gP��C��Lļf�au1='6�@�J�(&�O���1y�ڸc�g�`;�3lg�K��3�$�ډ�*���fg���xύe%iLQ�!h����q����}X&M�|f��,�w�������]'����uzN��@�`��D�@��^ˋ���K{�$ {\r �upo]�"L�EazN�M_Z8�h�6w�g ��=� d�]ٓ�4��fo�%��P]'&�sHtdO^ >@�|W[~{�o��\c�:1������7��z�����KP��(����wa�� 	��
܃g���=�&�H֩U ;��?���
`�I�<BQpO
$��ȋ
܃��OC$�� ������I�H�?H�o$cyY�{�x��%^$��^��! �|r5���� fN�$@_r�0w��/*pz�u��I_x�?X��B\�����<���r@9p�H*� ���߁��!ޣ��yp�����Gf�X�fb�_�W �m��R�I���.�H���V�l��G�� �=0����=6t^��}���t{�����<n[?�֧�N�7O7�ċW5�Z��C%�q�|�CWM�Z�=�R3z�CO\��; �� ۏX�y�C1wl��v	>|%��!`@_��
3���Pf((�X�wF�p� � �V��
�)����b�C���]2�L�&��a�ɰ�d#�D%�#}�.�9��S>K�ο�%�c�=������v��|D��� 0�/�p�=s$"E��0(�����^�{��0��o�������T��3�'.�p�/��(ndda1�:�����&&)�F��:��|�DB�0�o���3b�Ĭ_0���Ы%`��1�P|�����Y�&z��9���޼��
9t��wO����Qh(��"��=���V��=s$�K�%���F1�/�ٳ�U9� Idc���^Ez�<�E�D����I��8��S�S?���^�&jQ�ھ%�ڵ�u���h�w�{[�؂��c[�؂�,�`�E���ng�؂��U�}Hp�~�  �>�6DI{�2�!���(Cֹц���"d	�4�x�N�g�>Kh���*L����\�}���ïW�V�������ab���z�A��2��9���ä�{���e�?�~�+B�	!B������Dԡ������9��Lb�	P�*&�F�XX?啁Q��F�|L���_�=��������]�2��:�Tb���I��2�+&�D��2w��a��+s�;��B�5ì�1�w	�qe�r��9����#\�b�߃Rd>���_��zE�XD�E�XĆE�XćE�X$�E�Xd�E�XdE�IC:T��l��ԱL���H%>=>Z{�-ò�Ǧ��O��U�d��|Ғ���46t88������aYn��ˍ��k���a��G؆�G*QUE-t�ga�6!M����dK<���c��|���}�	�����?�}L��l�z��|����G�(���f�گ6�P���ۅ�R�0M��k�BKI���8K��������B�xF�PZ�Tׅ��j�Z�8��n��ա����6�UP�4�=~
_U�m�����V/�\�~��I�Eg��t����d��f��o�����z���ow���-��r��^(M��rn$Y(&��97��䎈Bj\��EȮ�ǥM�5�e�7�z�N�h��ђ�O�0��Z,5R��s���|A8�,�pfNke�#��C��la)!�S����2��| l�Vŧ�� ��h����P�%��+"��/QO��)���J��a}S� Wϩ`͌���?7:S^����S"�'&������Fin<�D����de=���F��胒���R�'��#d��h�Md	���.=�6�,>�aZ��8G$/e��e�J�Eܨ���Fx=@?�
�k}`P+%X��3�܆���O�������n�]������9��g�������?T���^�ek�����������ٛ�=�|(���ϫݪ|���?W[��Kb��n�����6ޥ�V�ڳ.?~rۿ���:�*=TH�~�Z@k]�R'|?�"�7�s˻ �YS�ʆ�Bgƍ�!���CP![T]��8.��iSmYX�,U*@�T�쫑F�@S4�Sh�OqM�M �c�h:|8C��H[���W�6|�V�3m��G;Z�F�`�ӂ~�p!B`����O����V[北!Gh��e
���>�=E�R��Ϧ�E�t�ϧEh���DAX�G�RR'
��R�ڮɠ�c�q,�>�*����F�C�B�Y�ł�9�{ �\г�L[M��b!�tС�,��P|!d[��eC�����U��!��&QO�Ky�0`Bu9Q/D���(Uo���z��N��<��gߴ��Zv����Y�Ø�xw`s>�Դ��:���&��^;�!h>�v���lPF�[�0X:|i��S�.ذ��y)q6�<���!o��Ѝ��^���ۿ��nM�,��l7�������p��i�$1aИ>�����݇4�U�\���L��u#�5��փ�
rr�JXڟ�1�����bpk�9���V�φ��<F�����i�B.v������D����m��p�_�$2����3)�ӋF���̓���	
כ��g}�k=cF�%��S4�=ϱ`�WdA�k?��f�?���/�q�� �}�X��W�7_}����~��gZv�󐰁��ǌ���t��a�4���R�s� !�,�e�!t��ژ��\��>r��_?�GBŃ�g���G���R1K�A�1��s�;R��`O���0RU�ԕ+\S�q�����
!Q֫��l@CN��#b����tP'�,��ǔ��T��@%v��N���;�&s���鵟r�fab>��vnB �SZ=V'�eD�0�
[y��0�_azِ��j��A.:�� �V�f����L���8��J� S���
aԈ-1��<z^r����p[&r%�g����3� L��0q���<";+�cGHsFZ��vcN%��J�$n�/�<>��M����Q��<��x����Q4gLD�����2"��C\����Y�VX�a�b�����v�q�ꃯ�9m۽������W���+�k��ݬ���w�7�f_7M|�w�������j�m��|�����EQ�������cN݂�ɨާ�j���Za�{�n�I�o�Ƃ�<c�}�K��qG��e�;�Z�3OT��bgc�v���/�f_d�;�}�	^��_�`����o������<�����I;^��x�^���B�Hn� 7:�v��y�"K0:�����d�n��z ;ڞ �+T�v@�=�灢�Ń��	���� �z��<ͱ<#�X> ��@bY�D� )5��S �'tj)27��!� �A����	p�7Q���B5���a�6�O�a/��N�v8�z<�u�| �"��B�\ ��H��4�����ue^ Ƞ^����ʷdI8@�P-ג%o뎓����W-�;������$|3���]>
��+�p�n�(��z��0�
ӫ��%��~=J�i�� �z�#�w�8LA��%qWBx
rW�w-⦇꺡c	
N	�jÙ�#����:>�
�^���#�`�W��������:��B�WF\�7�p�����h��X�]�:X�B�W�R�~5�z�^!W�I�;2"�d�6`�����Ʀ�{qS=J�8�{���z��������u�t�n������DަW��2k�M�����iɜ��C�+��:{#�-$��^5��4��C�ՠ��r�r�##m�;��K[ߘ�3G�Zj��d4���L�i�愇��ܾCe�Ǎ�#8u�.U�M�Ѻ���R��}�%�ol^
Q�c��=�B�\�m����[��Q��LDg�S_S���u��&�F��� �
�r��ůgo4���|�Zbԕ���V-��
��B�؝l��q�r�j��q�fW/�`	p�n|����:u��w�Z��_�Z���6z����R�T @n��9r��@�����]�;W�vC!m����m��@�ڡ���C���zIT��.נ^b
v����|�芳]W���<lm�/����No��V����ʰ�Tm�U��j�.k�F�V�pԫ�Ks�����; $��zx������v�v�74����|��[?��o6������\�̾�/PK   �-X����%a 3c /   images/26e5b11e-e137-4512-8967-7e228f6738e0.png��eX��5L��tH3 )!�]"�14�0tJ7H�-CK#-1tw��/���\����0�5y�眽�:k�'RUY�라�:<��q����z��8x���$\�(�5�;i	MO��6�4:+7�{�]r���lrwޝ�:q�D4�`��sL �~�����������%��F��"�n��n�(-��[�C����+����{�L��ת��e�K����V�@�wHtx𑟤�5�����[��{���_���R���C|���g4y�����I�!qX�7r�P*�?{����%؉��*�X�W�{�v$�h�%}�6P��,O�9/M�e+�% �t#%�xsӭO���ho��,-A�ɍ[M�v:�<:ne�2<%#}��V�g�X��ՙ
�&��m��|�`sD�;6'0uZ����8g����*[j�.)�L��NW`>�nJ�������ӛ�� k;;`�p���b�A�^ 3D��e�q�l��`��MNV��p�ܸ�����v��A���P�.7���������2j6VV�.�V��ﶭ� ��������rλT��KRv!�"q���ō�J�hJ�S���r�B/#����t:����'[���xu=��s+F\�=���.@�)�Qc
�s������'>ɭ[���KmGR�gW�6�(t;��kc8Jb��6xo����7���4���`�9v���	����| Q�w��<�#�$��O�_�u���"�G9z�2	�� �H�����7���������ė���~��;�?.Z�1D�0H�f�����:m � }���N�õ�k��Ǐ�Fc��Ot��]��¿����p���;UV��a�T͚y|�m-L��].��E�P���Lw�OD�|��ZY�X�xMz�aX�s|W,��S*�_|�����V��E�a����B��rl��A���2�͔g�) 8h�n�iڱ/���0����<}�����QW�'>%�S-�_*z1�[C��5�u�Ngy���-�� ��;��1�a�D�<��P����+m��?��v��8ԍ�.����S?-�L�[Ђr⍌�&�_�uBd��p_�b��U����l��:1�� �n��U.�ؤ@G�D�0-)����I�▥�v=�m���՟��k.�	djG/o�8��E��N6D�2�	!ބ'��cИ_�jB?�����oH���(����K`�� �7�[�O��Jk�Y_����Kʱ#���k<g��1%��?��	�JV�O�kt��n�?M��`��]��`�)���K�o�⎥� �����*ޗ}ZO)��+R�6�^�F�k��*l�|��K����IK���2���cg�{:]@\��pmX�ZX�PN��پwi�hVپ��-u2��|S�$�gvԗ��ȃ�cd��>�����������lIk�k���>T�P�����+���6��p��*݃�u�Da�}�@��H�a۰^{��MTz�����]+����2�O��9�ÐR�/�e�!�6���a��C6V �rqX�8�8�(�������x:��<��ve��: P�p���`�}M�I����ɓ��\�$V|fcR"�7埈b����3��ef����I|�Xa�E����?�ImMTc�M��Ѿ�/�Rke�5�J��&�CְR�02������_[��|ND�8 �C��h�O��ڟ���w^����QV޿�V�?5Gu�����Â���a���`ǹ8���P�8!B٧b��$��a�e��a7�~�<旚�5�G�c��=�b*���u���x����R9nZuE�f݅K6�.��a���Ӓ�9�PL.z`�
}'M�P��R8��h�c8�,r��a){N�aY��+�6�PIx���V�~Ҽ�y
{����T���+|3�ᢷ�.K�)��{B�Ý�˭�+)�j�5S��,C[�y�lr�ɲ;����yS�N�x`� �!�f�z7|��xǥ�k~��y�;GH[�$�"���0"HFt�J�h��X���ߪ����5e�)��s<T_�2��.	Jӑ@2�N���%\Q�O�V��H�>��K%7�9�E����[m7�#�Ћ|�w��G�	IoV����k�z�qs���jB��%��|�wa��;$��@'Ww��U�37y-H���� ג�Æ�MxX��E�.<��]S\�'�A�S�C�[5��,b$:pqږ�?r��31+r��F�������GV2���.���{ɶ�FdŧX��J��[ ���1�K�:��ɧ4e���t��
�7��sQw-VBW�t��\�0A@w �%� /}J� rD���bK���L���m�yG��G�|ې#akͧ*���E!B�;S��X�7���!�'mb5�>���-_��^�j��n�R��`>7��'�v�[N�l:��E��d�(�#m��o��t��R=�C��vg����]}����l�ʅ��Af��U4x���F��L�-,f14�w$�ۊ�S�����n�N6����K��ɖ�O��ƾP�*��Sk5C�>��덹�)��w�9���L�E�X-"���f=��4��@���,\$�)�H��L����rt�uZ��Էo�h7>&����}'���1q5�1�o�� �A�Y!�w7w�+�;��U]L�ۚ��7q|�	1�nqMZ#�I��D�o�� ������r�����a�Q}Ss��G��_<�[3=��+g2�w�E,���R����9<�����=���j?X�~�Tqn)|�a#�����lX�vi\T1��#O��t}��5�)�7��������S?l�O~/���Oq̆%%�z�_������b11����!��s/Ī|���궗d|�4`9��O���W���1�I^��h� �	�r�~w?��4Թ�v��,W�Ӷ��ӓ���x��bπ{x���Cر���%�g�_Q��n�Z�`��J����x1tI`tX����B��d���ⱽ��A�x��/�Jxb5OD�]���>[Kݏ�����w��>����>+�B��G�|�L�'I���Z�� �&�cQw�����.}��Rt��&������"�Ѓ��H]4�X��I�
 �Φo����y^\���v�׈����o6�*mW槾� �?��?�Qh��Wfu�}e�ض�/&vxڇvD�a�E���U��\�6�aDA��!�l��Mk(�)E�.�7�s<9#���a�o���7.�;{6n�P»�m
���t�8c6O�7;L�R��B�o~C�!�1gP��]Zo���2".�jc�6�ga���:����9F�頲��y��:Tר>d1��/�4���"� �mr���.��幑�v"��2���������0lT�+4�_�ӄ�x=W�Ƽ_�>n���xW����%�?�EEH�c�Z��Ǧ%��P�@\hR/�+M��&�a����I���&<���>��o���^�Z�\ӗk-�V���<O��B��'��q�d��a��xI=�m\���I��M.��[�.���W}N��$�I{+�;^�`�3¾��6�����O����k�G��s��w�r:�Ƿ����$�R���������H��k����a�.��1�$�ڔFG���V�l-��o�'-;����j��ԉ#"��Q=+S�/��|�vm���U-�ه�g���KYg#����Ks��/RѾ�lsӁ��޿&f�SNs���e�5~�]� ��]�5���Z�k���z|ZZZ��=���wad���\�3�C��¤g6�`�z�z9K+j�$���3�!c�z

%������z���Њux���!�:��3��D��J�/2VZߋ�"���Y���T-Ԛ��$r!���|/kjZ�;Hp�7p_����r��
�\~���,�y/��-f���k$���]��3����ʊ㒪aA��P'��m�7���C^��U��b}�!f	�ӗp�ЕH�*z[[��&��9N�>����^3�E�+Bzi�l�;^�Ǩ���r7��r�/Qc�w�3�7j_��`�js���xt/�l9w�b��S��9p����M<���/r�U���Ӯ\I"����W��y���BB-�/�o.L��t2�ݏ��FȠ>j�M���Ԅk�'��]2b��:#J�w��i�L�9vhO�}Gm��ɡ��fA�϶�0��?���aˮz5S��Z��^0��!tI�k`��������S��gu���HTj�7ݦ���l1�A�"-b
������E�NZUb��#x S�d*_v�**H^Z��2���U��gdl�e�^8���ߔEF�!��9�/�N���=��K������7�:���"�j�����Ҫ�8o>ΓUI�վ�R����99F�X3�3r^���V �8���>q�����f��r�������{ �x��9�h����O��8:���=���������&`U#���&��hY���M�y.#���E���F��[c�^B�b�x  *s}��:T����ݑ9��c�h�3о¨�9�!��ȓ̎�}��w~VkC-�F�	���t�f��7���>_�����n����>i����EM�{��y��8`Ք7v�D���(��"���~<�bŉ�����n���vco'��d��m�u�t4Un��2�C[nƋX�=�e6;��\�q���u�����1�l���:�ݱ)�YP`�W�`��a`E�#�����Q)-�/�}�����n�(}O%Z�f2pёq_"ϾP΋�*������Z(Ӫ?��rJ�W CD�r����k׆�l~�7�L����ߣ�	ܥ��n�]n&�x,^�����������xt�b!B�u���-��o�¤�_�e�w�8K�� ��E��}�{f����8��L�Kb�d�y�cx�K���}�Xey��KD���z6�!�cS��{:���$�Bc��L�Ǭk��u�}�1
����6����.����"��l�[�_{�3X2��7����y���Q����P�ɢ��m�2]���m/'�7/"4����A�G�� �σ��@[J�tR�����H�E8&��D�����E&uM�7�ͼq��h�#��=n\?V(������%!���a--	=e��ӓ�!8Xx'�(�ok�،+����[su"8h��P֦��L��A�{��a�����OU��}3��%�4�癙��{���;�n_�$������f`^�1�j�!w/BZr��m��"#o� �YF��E����u�ϗ��w�����i����K[~���\h���l�΄r�W�n��:�`�+��
��*����iYk�W���0����=s��Vb�?.�|6t��Mg��7YB'�쏻�ݦߐ�3Ȝ���v��Ü0-�g�cccul�d��`�Bǝ]��.7o��y*�lQ{�-�q!r���2�ԡ.%"X�)<6�kY��]A���R��ׇ���2j�^K��"���r�_�T�#/������<�N|V�k7���/]7�X�i�?�b��M�/�o��0q��:
�@����Y^�G�~�f	**�]���v#�1����\	���C��U.]K28Qm�J֣��[�|�T�,d��� ���YBti��E��ǫ�g��qp��K�g����Bo>�H�����^��-Q�@M9����y�g8=�T��Ft8�,i߳Q�3=�*�]_��¨R�] ��t��ɜ����aqޯ���K��0�Z<Bg*�5��d�51�_�F�g�>I3 p����`�b�����=���7��ǩVє�s�*d1L��F�p�H�ƠR�c��PPHp���a@x2z��U��胵�����/�c<�zTr}����<5s<r�x�[|�&��O�����	�;���:�'�����(^��/�ּ�k=��$}e���b�ve��3�^���o{�+S޿���������)(�� �ʃY���X��c�s�����G�� )4.hz_bY�!Ԅb}A3,�L~����J�o��bW`���:A�?��쪫T��]�rF���;U6�@�\���gG1�1��%߆�[�&��%�-�-D�hq,W����&��u �=���՟�!���{)�ն��.xp�k�"�(��t�d����&o��6�.��k;���(�b�\'l��f9ND~��^"� �o�)ް_�<v>c竳IB�z�i�^����'i,������$i�F��`�N�ԊRNѯ�g�=	��/lB�i��LW{�sX��K�4�Pev�4צ�E�*;�{�_ۺW�'�@du����d�J^�{�<|Y���4�<>L��1M�}��^�^��һL�1��ұ�:s�������2ds��P7k�\��p	zй5C~񀟗�r� fV��^E N"N@b�w�r���i��j�*V��7�A�6H����'-�8�K�������q yt!��,c�����c�=����2� �F��F���̉Oe�>/����4�[�g�X2�?[��K��h����Ss�c��Vc�8t�x}|��W=��Bt�b���4qm�O��3}��n~��\����u[Ha%�=���
 �3	2l5�c���'r`&�Mc��tZ�;<��E.�O8�p8	HȔy`@��m��9�(�b�mN�A�~����u� �^V�ě���::{*n0��a�*�qY�;?�%��^m>�_�ܜ<��EZI�N�ԩ�T�4���?�	�¹�^ ƪ]]�V9�x���� x����N���vB��t�2p,����	�n*>� ��Pyg�6�sZ�`�ؚŎZ�=�&,ߋ��Z*\�������ڳJ�t����X$D�-\�0߈���\1���3�klX)x��B�~��W��▤Aa�h��%�@�`�O�ߤ�3Gu���mp$���,e�����9
L�V/P ������H��,/�1C�g;�V¯DF7_ńx}��wy0��v�aB��x�ķ�h���I�[WS�j-�^�d��D�=NC��
�-��<}.k���`��x���*�[�7�"��ȫSp�����d��9�4�8�R����פ�7-�N�CH��!��X)Y���<_��B#n4\WPQ�݊�W�\�����QT R���N�C��L���Q�gv�#�?_Xi��w{ѥ��d�ƕ<��Ÿ�oOv������!���C���5����Q�m�yK$�u��oK$��<֫~�-ۿ#�}����TC��.�ʽ¸%]�(Gk�U����pJ���!Q+�>\�*��l���� BYPJ
f%��u��2Tmy���4�I�E������A�ÆP�@ b��h�	L�\��~�0�}�BL�O�d�'qꤷ3#[�~�����F�Z8�x�ii�ǃ��.��x�Y3�ƣ#�25��>}�W�^sJ{�
d+Я�4��1������ä3sF���E9�0�hW��LP�z3����@_e��k��:���`Q��t0B��ͮ�](p�E`$x�l��K���C36�V��3��nӝ���,�m6���/������������b�m������²8��5W��¤O�[�
�@&��[�!p��J��x\w�宯�a-M�>��],˕�=���v���uBv����}�lʑ�x�c�WÜ�����e��نл����B����+�����X���� w�|�@���P�J=l&���)��� ]r\45�_:FRﾳ`z��v�d�F4�O��|�����;�b0�4 ���H
���8��E`�;���k,��-g׮�NCHƋij��3��nՍ�-�F
�������fٞi\'O��л�nQ���h����^ �tR2�;yƁ=��3���a99تN/,�b���9%}Z�YM
J�zc��g+2gٔ��6��B�ك�e{�"�'��T�&#�*�a[��UY�/�V^���h'��::0'4�l�[�|ݹ��]\��M)��+ �c!:977� �b!��E�i'a�qwK�m��\g�$
W�x\�~\�	ǡ�!��a2�'�iB�s!�(�����kۿ�~6����F%�� �����lWRo�Q��e��W��]j<���z�C��(v�&5���<B�[�� ]	O� �흝�o�>;�B��#�W)\6�DMꯝ�F�*۲#}�����}^D���y82�������<�M���'��\�S,�^Ϣ��0	�O�*������^]x|����Iwi�G:R�<TM ć�W%V�lA+����x��.ّ�	�t�����⤓*�8��!�v�*�1Ne� ���ֽz�:���g	Nh	�/'9���	�?�@�8i�钢9V��m���Ȉ�fp]4[k����Y��gCk��������k,��.�a�Zī��O�Z�7�g��T˵���O����0㝷�Pc��)n,o��q�CZh2[�~�թ�k�/E��Y�6w-W�鬦�_�
Ü���H���<O.�>������p	�z�_�6x`�JJP����x\y\]�|H.f]��{V��x�I��z8v�ϯ��Bn�O<Oǝ�$�1��ڏ���!�Q�l`$�Q�"�$?�؁ء��߰�$Ir2�Qk�x/..L,�_��Xr�����p�ph�Aqp�@�	��c)�cg )�iH+�m�n$W�c�W�R���d��� �}z;}䑩r�Vl���#��AX�Oہ̟>������ٝ��R�lij	�ÅFS� b�Y���C���|�(�4֤�Q,�
�d�"W�qTbq�a�v˭��t��z9���f��؎��#��D�s�<8Ҏ_u�W�☈ޓ�('��<�F̔=�v�m��`}zH��j�&Ȭډ7�ͺ.�M�'�,�����Q��:�p�x���U��B��(�pbςϪU#�P�RC��.Ў�� E�2�rs�ٞ��?ch�͎����d��G0�������
^y�����x�Y̘k���H��_c%��U�\EWnd�cJ']ϙk�Y�ʟb�/��SO���5��C�M188��\`�<�wS@�"f����juA���6(���htv|�sʳ�]ߖF!��Q��Y���Y�q~u�>��`5)�1W�^�J�Z�;&�r>>����td�p�ǭ0�Eg� c쌎���� �R��L�������6�YEz�kaHG�ï��۳����7>���Y�PfKC�0T�E��<�K��X�<x�*��M������h���*��UY�f^O�W�̰o�F�LC(P%�����]�%�Ӌ�uv��ZMQ��lq%q�53�4KG���^�J��xK���>N=)��2����/rl�/B�}LL>E�O�j�^��F�������Ē���< �����A�`]���?��֊=^�r��A6�p��	)����9������9ɔ� F^����rv܀_ꭟͨJ�M��!��m����R��E���d��T�lX��t�=L��ѽa+��P������y�(:ԥ�v\���Z$Z����D})�Őᵼ�=��>��d����E����1���n�\��M}�D�˾T�������D�㣿���hL||�Rh^e��W`y���ԟ��Ѫ�&<�ŧ���d�����"@��MLkxҒ��)��~��n���A9s�}8茻��Oz::�\�!���������0�Tt N���ۑ{�}}�����0�ff�/+o3�%�bd;ƌSfsvT�d��.3I�*��;�h�_�H�E���wIV��X�p�~KQ�}��7^N���ž��������9���B���OZ��ǹC�X�6���hl���#��%�U*�||iid��\M�[�m�o;����@�	0���e��ݵ(#n��D�JY�WT�m0�`/�d��م�>�}zOA�Y\�̓�,���Ն���p��#���0�y�F����1���ގ<#������T[@���V�S�~g[R҆O�J�2�P�g�)E%��	"��q逄���g<���u#'R_�����-�jס���	����yiǽ��Z֦������ �"f�9�z�}K6�����S�~���%����B7����ڪ�JC�b�ʣQ�b��$�gAy-"[~!z��7�V`#�+d�*bn�+JD7)���bu��}t*����O7�G�<HM!��y?����q�.C��HkI�Z9��`o����o6Il䅆�nQP�\$�x�A�:SP�w���L�~�ęS��)_��{�q���'"����K(��5���1�e�g��T�����eY��6٨B�������`���ʆ#��6s�
� ~&Z��/3nC�Fm���	2�`��@�q]�T�C����B5��qZ�+M�m��e=��$�����eHi��� ���5˲L��T���Q�f�`������cU���_7.��j�Xzs^�Bq���kjΛ�!XKL�!K�5]���Q@{�%�f4NDå��PR����h޿8��:�5>�c�VYH.+��;�y�@x�����Ã��d�ܦ���&�n豓�"-L0Z�R�p��q����}�|��쓽���*��0�jX�/���?Sm��&��+���f�N�����d+��2�T7��n�ۈ2� �C6�#�B� ��$�*u&�%��	o-4�P�Z�8��T�"&]bm���{[G��f"��4R����X����	=�m?��ݏ��ڳ=��8
�4 i��|��������4$'u5��wH����r;��>�w��U2�9sدɊp1�T�>�B���t�L��E�4S���5gw��>�#��A�[ι哫N�������c���h���p{k����ۗ��+}�h��W@W��NQc��G��d���3�]3#�ۊ��ժ�q��UK�~7��M2�dc.v�ܠ,:=|r1p�	N��aPw�dM� l����-q:�׽^e
l�(�#[����� M�^A!�έ6�w۩ח�V�M8%��Krq*O��`9�ü��z[b^��(_ܽ+^nnY���3�����>��0�['z�ה^�w*�������zoRZ�ye�}�_��w��|��.���&�_����.�y<]�P���`�$�"���׹f/2�wʧ��ĳ��"��9L2�n����E�=��.'W\��8��i�~w��ĢX	Ť/��A�,��g2}��a�d�g�ىr�Vl����V7��w�x�e���.?��d�f��2�[,�:�a�}�]�i��H���^ϓ�j�Ѕ�	x�H������J��0��Ll�N�v��M�_^���&O����vZ׍��UW�%R�*��2.��i'^[Ii�c�]Adw�����L���:|��&�7���ߛ�JW�\�+�K݆L���k� ��՝�]��n�f=� ]�.0���nJ�X_د���|`�+�l ��e�����Y�O[)�a�T˒���`��K�,s�\)�����F�ۢ�U5v`���3ƥ�3�G�8�SG�֖]��o\Q�?��M=?(u�����t�{�ov��~iwo�l5�r��4� ���3��W�U(oa��������������vQ��|�k�/61��]˽�Vֺ��P���v5d��� �|K�W&�
k^�t���u��_9�X�L�Ew� ;J�]�+|K��,���ދD��3��t)�t��#`݈�I1�2��|viڱ�U��G��Y�GU�.�mܧt8�NG��AN�>������S�[_�����-�'��|V`l�������7��Ĥ�r�^���j�돮#����{mv���B�3����,�ɑ���vrO�HE7xO�����P
#|584�+@����8@��얾1�޿����`дm����1�n�GD��74�����K1� ?<�:f~�uޱ�ݜ D�V�-�3��Q��2����oD� ��f=�J��kEO��e Q0)�%��1*ô E<Põʹ�+to�~U|G��NuK����h!mhv`��(���U�;���[#^8"R��-'.�S�z�	�h���X��"�^�ը\o1[����
ev���V�r���'a#Ӊ��;]+�do/R�}�$�K»m�����?�{���>�l�3���N�bϕ��p�8j�����p�z���(J��$��?�F��N����E�G�%8f}�3�z�+��a���!n��혊v������8���`�YP�B�����f���.���BQAC��Xg��	�1+���]@x�9g����y�A����c	ߑ6���>ew�/�����EED";.Gv��7H�#W#���!33+n_����V$��d�Ԓ9�Z'�����P������̣�>�r/��xÂ����>�H
��7�Q�P=�=4�4{�n�HeT�9��wEr���H(���}��*su9>�$��B `Z`���k�-sX�@?<����Cv���Y��h�)�r���E�h�7��0i�̇��_��wtfE����k/.}��7:��$i�RcJ��4A}��V�w�oh�oI:4�Y�c�� [e�ٟx��T|�,�Fr���UU�2�y԰V�&A��L0�r����)����]�Z�qKىٗ^� ��EByNcT�
��K��rp��=��t��S�r)��)9ʾ��K���d$Ɖ�Z�Q`s�&Hs�x��D�Y�~�k��e`:��5���~t�9>�+����QŌf-���������z�@U���4�^<�F�>��9�*3�/�[O��ӓyC$UV��w���˗��\�^�tGj/�R!��(�[g������+R��,|q��tt��]�t��1�蚫/�bHvD���N�H�F,Gv}����$��X��pTK��k6�[������o�4�����)�F��is��X9ܬ-]?V���]��D��ɥ!����m��f�J�w&���Ч��d��4��n,�,]��:��C�VN�p�2hxJ�$�����v���W�R�iݧh-��h��@�d�Wa��Aw�o���B��s�@ ����\d���X��~5��V�]B�`�+��*r�HiL��=~�h���@�%����:�+$:�[��U\`(�ū�f���=����u��a	g�#Օ�ۯ�w,��Q����jАBpj#�..֛���f�����]:�n 6_����лh�E�'���ӽ����1s�Ha��y��pV[݅���5�>�nU���nk�?����̪UEKgÉ��XX��ٜ}�� �Y�GG����u��Ѩ̘Q¦m�>ܬ-�N�ҩ*I�'�D)~t�*l-ة1x~eت�o����b{�Q�d/>�(g��ay�lq^�&Q�
�|�h�q��B�3ӆ����:�TE	a����'�ӆG�MOd�^���i�.������1���CI.�y""�[����l�������"�z^ݺAr-���^�^ F3A��
���A��`���.?�V�`f�ő�F�4��܊y�a ��]��a�>���RQr@���{r �r����	1W�,�9��HR4�����[��;�b��,����C���X�!��A��g}�.)��W)�J]~Q��Tz���>Bv���I�~��9�\ �~����:�c+.�y<Vb�����r�nɷߣ *1}�,���"I�L�ygɍ���9��W�u���Sm���Y}�% �:!p2�nR����c��:D}����H���i�N@3Ey��ht��\!]�I��QL���1�lb�o�DSC_J��Q�S�`��i�S��A����B鳦EzK��Y5�Ea�� �)%���1�V݇{/�ONpC�uX|�r��E����hr��yr���&iҾL堲��5]�0�.��B�W3��+CL�TP7ok�$�±��,4>���<��C3»k��E3x||�����M�8c��Ⱦ����$wRE��XII^FF����&�'� � ���J�d�\;���1��<��k"-��HFs�}#���/�s�O�eM�4^{T�}H��N`!�FpRO���R�Do�;
�J���ь5�&����$� (�M�f��|��:�{��wg�g�6!���ʒ�*3#�[i���{|�;��umj�ZN�M	)�%.Iig䰡��GR�BO($� �l���EL�J�t���m�%+��������Rw_K���k,������A�	�_�#��?��K&XfHe�F�V�0}J[�T��К����q��
��ۙ�Wb5IFh��+�B8ʵ���B��&nuP<L^L�V�PP�$�����骐����g2�[��:L:Fk�ϯ�!G�<1� @p1�9��즕|s���m�p�9��o�^Nغ�DͿ/��N'���Q��_x��v�.`߳Lp4��=�Ƃ�P�~w����O�Ĭl@{����t�X� e4����������u'�l��&f?�_����o���<�ů8--�:���=�]���T��c|83e2�aPi�	�yi~F�rawrK���ֵ�O��kH��CD����<�Pƛy��'i0�%Gy���Ŗ�|z�Hz��Ì�"n�.�d�,o�&�.y��p�>Z�(;��1���=	�^�CW��ũB��:��W��^�b�CK2Q����f8M�q�SF�h����Ē�b30̾>�`�yQ�p�-K�����X�MU��bO;;;E�s��Ss��67�$?^�N�M��լqUĥG�B�`���;��0o��x	�5���Ʌ����������D�:���o?���"���r^�"��6�XYYA*�Z��c#�X"`7 AAA��= [�x�rlx���^��<A!������`���O�Go������lE��r���Ukz>������&�COٯ�b-�㸔�������e�j�@T��)��
XZ���{����(����~��.t���iɉ]z���6�+��=�TB��N����g���J(�T�8��@l�4��eu q��f����Z��i���>�S�h��e�;��2���K��l��^FIzzK��)&Eee�kϪ�9q�"�o�[Z��t	l�ՁLi�AO�J�XO���T�@�3oq1���+�h<����"�.���~.�as�Q/�;⥣4'��>���KQ	`..ik}��w/nj����}���}\��w����k7;@������}��`7��'�[�Ϡ��[���(��[�+n>>j�	l���b���@��kbt O[͸�(g�G�Ǣ�����]n����jO�w~x`�KMw�:=g{�����7��n-�9ܑ��fe��?�0�.�}���2�N�9���Uh����y'�&@�!�2�����[��q�S�[�~md\}ITd���l��L����Ȃn����%���w��p�����1��KH�h���H:��||�n�ց���3����`�"�Л�3��z��C}w����ש����a����,�(߱>�����h@�@b���ǃ��P�,�mz�����f U���S� �s)�!�fu�{u๽�0�ma>v��[
D#ϐ�p0S)%��"�W�HH{6%o� �6Z�<mJQs �w懅�|�@�v:���;�I^�fO��>0��P���z�&�Z�%-8��"��굲�a�� 9!Ș�E�f��ȉ��C�c�O$G��p����0�~�Yh�r�K�/��X��y&Q|,�q>�!�9�S�C������[�ɏ��讽� ���ݏ>�1����$���Wǝk�5�F��©���::��F�/��*���	LY��OgTV�!��=&���\"��ۿ�8Oc����s�b���au\L`��v��pJ4:Aް�LJ�:�Qk5va��I����kj�zgΞ�#?�{g�����ND�������5����3Cw�	��NI��HE��b>����۫�Z�urnR�
�"U�*�n*I�$н�����o�$%OAж&�j�ܼ���l"�^ G&�ƃ�˷��D�"rq�����\m)G�R������%,������~ �/z�x�["վ>ﳘ����|ܜ�>��M�Y"=[mZ��w�$q��6����[N1�
��~�ᇇ����E���7=���-�o��cx�3�ߤt._�J�3�!��&�� �.���|�%���[h��	.���Bܕgqܡ����"~�5��ǉ��2�$B�����<�i,��W�F/��\�^5�8���[T��.I�לR�҅D-�E���-s�-rӃ��S���	֒��R�"�-t�V�J\g�|M]��ke����Q��#��+]�~��u�c���"U��M�"�-Ř�j��9�靄J��^�L�B	���1pzKY�,Hy�������P�Q��Zz;x��W�*��^
�(����+s.��G����3���B���dp�JL2��[�����z�$d%�b�+�ʞK�<#��8?%���0��v��g�6�6��C@ޅ�M�X��	����-�}��)-��Y3Y���
g�FD(����I~��U��NH����8ª��=����1�Lq0��(Np��݃�;w���AwwY�uqw_���wN�[�������#yf�z�xh�$���E|�̜���a7'8ǆWDYSŊ~�%�3ud���su+�c��k�
�������$n�R/8��t��N �R����@���A�M��"G����D����N���k�g�O��k8��5F�����-]������ OO�9�B.'��J1b⭐��e������[�͓�
�������6/''��+|UF��<PR���E���^�y1��o�_9�&$����s�K}�a-j�%�fհ�Z�Y��ֈH�wd�j�_߿�e�z���|���FzZEz�A1�}vN�[�'��e��e0pA&���շSw-�M�0�i�cG�}L�X�pJ@��3��$����YG�*S?���ۼ��RJf�-OO��^�ߦw���d�q�?Y�U�|��%����6"�ٔsy������}���z���C��7s��s#׳�0��J��[�L�=�?��89y�@?�o�L�~��edHI5=R��*��]I&MD>3�+�=xt��tY�HCp�n[5ۚa�F|��t��5�&��>��1��d���E�l8�֛(C����KY��ʍ�ԙ���$���"�`۴��?�M" �{>��kz�`�х6�(��ҋl�"J�/9P��W���q�����B8��p��_��sHLE���*������m���\��S���CG�T��v��~��C��z��Y�R�Ƶ�KV����ۢB���h�,�k/$G�	���6�Z�Tt^����B�=�m[uz(�NX�� %iE8B����d��������G�eko�Y�ϒ�����#×= Ͻ���"'��U������7�����Co�õ�E���S�/[��ſC؂��\��c��|�\S5y����D;��2tXH��BۋLv��t�Sԝ��繥�V?A�����0����-�W��v#;�M\l��茐��%��r�o-���ކ�X7i�TT�|_�6�
9w)u���]��^W��,���4�,i�X�����E�� ����;��SPW$GO?���ozk)�\���H)��,i��;oJL����*�g���ủ2��-ҴR�����2�z�e��Z@)������V�H�!<�g�
�B�l���[�L�����^
�b�ؿQ�5��;�}I�����i7."gH�?����ׅU��1�o���?���!���~Öx��_
�_EiSY#�J&t��R�8��l���-�|������}���>@�	��/�/�B���pbn�8����T�s��x����1>!��JL۵'�1�5�Bd���!m2��G�+�{E�����|�P����^��0�v��W���=?�1QU&���ܨ�6M�^��?��6�dʐj�\R&xJrs�@��W�� ʇ����i���6
c���_�m�>�6;��\�F����Ѳ�1]�������mgF�q��<�{�'�U�>��������\m����U~��PWU����L� eF�C�;e�������пșb��Z9��q�e���S���K��{K����Ƀ~�o�w-[��+�퍡�O��
㋃�H>�Ҭ�φ@a�B7H���7մa��;?=�y?�2�1�$m�+O~]� :0�^/��.pJ�?2R�3�m��>T�D�G��+��cq��U��jd�p����Y0���J��`�d�p��Z��*Fs��y�x?�=�z��NeSA�O��_��p�q@8��0ȸ�ˍ���I݁Cq`Ҿ�h�s%��;0��f����p��2᷑�&�$�R�0��l��/��w��]��Cc�͏ѷ"3���/
��5�i/��+]�u<+�`aa���~)�.y�O�ݿ����Q62�/d�@���\b���I��i�{~����?�؏Ҙ��39ع�����7��*���S?ڻ�r�~�I�,T��@��-j�ғ����l�' �)���x;���)D"�묫�]��I�0���|���_�T%��2��Z!'?�X��K���_�V0�tDv��%��]�Yf�?ď�`Z^��ޅ���L5U�>dTx�"݇����Trq��a��5T>����KT��l��O��ͽ	��K�;��>��[�vyؑ��<گ�l����pG�-���e�c����M/,D���+��-r��4.�f`�?���$E�q�m��kM����1&[�qX]J2�7���a��y���y�Bs{�,�/A����<�6���l
�,U�^�f��b��9:>�%~e��l���3F��a�1�buUO��.&���z�0dB��� ��U;�::�������5�ԢL�-�4�u����.J/W��ШJM|ИFbN�c�R�R'�L(�50~J������R�P��6��sX��7�-���g�Lu�
�H��syQIFF� ��r��C��29�_���	�.6w�7�(t'����~��Q�V�o.0�,�O�1�ORU��먉�4��\6ݼh���������y�0��-n�Y��F�\NY�$�+^f?�4�B��a��u�BrG�
��k}������A����/m�Ă���c�N�����#��ɥ��|�c5�?b�4D�^F�@��|�q��,�oT����=S���������(Qf������ac��W��������=qT��V������O?����m �H>�踂ԡ�X��2����y"��5&.�<+}�P�;[W��8Ϊ�XE�(��q���,S��V���2ir��M����h��W�+R��,��9�~��c��y�!)H��S+/�"iB$>�	#vc��|~~�_cHjsw/��@�����5����h�Y��,�o�f|zHTN��0}U��/W��[�Pri��} �g١�^�������9l�O���pQ&��[�2�PZ�hUJ����b�sV�αR��E~W��9&����T(�j+�gH삣$�r���i0��x��*D��s4 ,싟w؇C�AS���Ņ#���
@f�.S�����!�9�9��Q~�r�'��� ��PA%V���\�6��4�Tj�rIq<~On�E|�487�t�`�A��-hi~>P�|��8��>A�CĨ���O�h���e����[IذQf�����q���!��� %�4�<o��d��t�I��#�%������n}��0G�}�d���.%�����y��r��\��mzljlc��_.\(��a��4f��2j�����)Z���Iy��ʤ=[1I�ʽ��4��	�6f7w$��x�q������oM,qc�9�����)(0B�@4C���@�m�����o��\���s���(�Y�^`	�c���t��-B
;l�vs�]�[�@M���c�
zg\5[���f)�
���_۰���F�d��[��=w�dϾ�O�yn�"��@2*��^ѿ�u��y#��!!��-Ejy�ǟj����Y��T)�3{*�?��@&KG��۰�o�ǵj�׳q�j�Է���ۅ� ����i��ѓ-Zկ���I��37Ǯf�O�� KK:��oΚU�&�[++�^�ׯ������������q#!.�-M�U����8g�)�ك�i%��%���w��i��-^�u��*.����s�q��E��_o�SNR�[fQXzG��2M�OҴ�������{V]'�t���(���/N.����F�����Ԃ5����!X)H���p99�V;6^�����<A͌Ucp�Y�~�k*��4jv2v� s��yȍ��p�p����H�e͍�)����>nn5'����y�F�����m����ٺ�!ϓf5N��V[�YĄ�����L;��9�[�P�5�W��a�Z�m�x��<����k�'f3S1h46��bM^]�Z��.8�)W�V_�1�Tl���I������Q $ް&�����U�<H�u�k����u��i�}��fy�l�z#|3^�7vs25���*�W�M����.�|41b�7���>y�z�����~>{o���kxq^����4U-U1VH6i��#� J�T�`%�l����|=�Kc�ND�/fi��0y�7a�R�"�/b�rx���<To%��?)�d;��$����gP%Vh�_���fqh�t6���2�"�^_�-�X?�?�;���lk�6�+K..�#)�z�%�PYve�O��y}o&Z� =��{=7��Rc����fY�)@᫝>���rU��"��|��<B��֏ڝ����Ɨ�`�����o�GJ��4lN�������眵��a!�Ɓp|����E��:~m�b�9��t4�0yf��&E7��6{W�g�ⷀj�2M�1=\Ī��.���H���x��A]�ptP���6��$��%����WǑ���V�*���~��y�n�L6���!�����~W��&_8f�ӫ�J�#��/����_�J����h�V�����ٺ�WI�$����H黬^��/��d�-JL>4Ӈ���R8���U���.h~��A��TJ��?��N�N��Y�,18i�Jk-.n�wt�<��*S9��Yh�K)��k��h�:M13�AS�|�������}7��F9�e�q:�C'�JG�xg���8� ��l!��(�$3�\2���l�;��dN,J6� ��W��� 	MM��-Q��:�cW��vw���{�~Ż�ұJ�c�����Q�����{{��ֻQ����u�̪�'���Le926��o�XG�lw�)i1��K ,�K'M�>��h�z�d��wr���!Q%V�u��!\������o�	��b��R����Q�&=�艅�(�Uƪ�>���n0��Ց�is\��W�G/7���R~�y��n��jY�A/��	�g�bMlRM�)�~��z�%Ʈ��@M}rƧF���<��#�����թ�f���������)�y�T3�8JN��?��^Y?}{��ך�<�  ��I`��͎�FͶ���3��3nb�����O���0ɸک^�� �Ռ���9]���k�
Mz�!Y�>�k�a������˧n. tq2��w�j��L%������kn�e�NK�>>����7�S�vkr����Pp�g���`�A_�n�:�d�x�M��!T�!��/:��n��a������y��M+-z/i��Y\���d�*1�[���T�����"5�x����f���i�:%,{��Cu�%��^��˟�q�0y_Y��N�
���|N6�j��Xwk�[~�����uC4p��$�q��Va����c��]���6�����'�!A�*g����.��4.0���C�8��A�3��~AB�������L�F�q��#�a>:n�ڻ�:�d���g����nbF�{7��(���_���m��r^+��ο~:@���1%˟����t�1k�X/��N�I�?���En��>�:a!v�ݷ&��u�����a�Η�S������o??�z��Ƶ�k�<��s�a�s��Z0#�z�a���k��Ff�/_��w����i�ۄ<-�JW��.M"��&uR`�A�X�\��A1��\t�{��^J�0ע-	m��ŝ��U�����T�O��*�{$`��?CP��+�Yخ�Č����':8��U���1�m'���@;�8w���c�06�(���
l|��ꐕW�!�3i��y��H�_�w���*cB4����cl̢�����V��p��=�5���rE�/����$,M��\����a�.�F^L;B�O2@��>+�k�DN�e�1�?k���/�4wǫ� ۹���ڗ�a���D���k�cb4����S<:n���DY%zLe�#ժ�,�l��Of���}a28�3��P5�%���Q���M_�I�nGI���8ja!-��ڟ<�P�q.>������%㻃�Ѓ��K<�Y�b�R��cy���l�!f�,��.^=��#�88F���n�Ш�-+�l3:���lӔ��P�YQ\n]y���P�h����h���е�[�
W]�YPlx2oP��X��.o���&���2��@Ύ�4�tT.�i±!�ǿV$ӿ��b���eh�\��|��^*Z\��f����k����g�h�����X��&��4�\����f��7r�6D�)�'+�n���A{��rM���F�c�I��/�|�����^���JM��oO���=aa2E>r�����RR�i��	0)���|�xW���S�&��Ӑ:�as{ז�I!	i�F�-̳����A�[7u2�#G���.uwe��l)��9	}�+t��
[�YZ�ӯ�<��Ȑ'�<K��P�cN��c�p�����O;����%ũ���;�s���,�����i^������C���]��0�r�rã$;/�0�7���/�7S�W�@ηF�e�8�\����B�x����L���e]Z@�]���C��/Q������'n�e�-���&��t�ꀅn|Q�G/k���V����qj�si����fZ�쯾�c8H|S]�t뻭4�B��n�k}��[Ҡ&7{G-�4P�V��c?cYh�7�M(�h�]�Å���σl������A�%/��L�8���8ěͺ�QA��ux/�=��HK_���D.�B��~�+B~�h���;���|Iy���bm�8���[Ri�ՅIS�|�%у����^�$��}�� �:��
���l�?�=[�$�YH(�d�\~~<�~�� Aݷ�%!@�� ��]����������r�xD��(��3I�~~wWq� K����mw���NQ/�s�`oo�õ,�spDVO�Bn�|��N�ld��y#��;�u`}_�\��#b��
+\߱�,�{U�[�8W��:I廘D/��X�p\�8����5'd�
�?VPϓ��B��RiQϧ�A��h)�����u�a��E�_7|�;��a�����4�I�%�֓ɻ�ť��?�σ�*���Ҥ�k�]Lu�K���?G���v@�tz��y�?�s�A7�A�ԏIr�6�M�e�+���x�8W/a@V�V�*���d`R�{�*�
�g��Z�'ՙ���"�3xE���|�;�Vgx7Y)L��yU���@L��S�^��˘٧�^Ju�F8��tb�3۱%C�?�f�J|4�}^b��$�/��_�KK��=AH^7��y�%
*�g^e?SR��GQ�n�_T�j��<�.�纆��(�ѷ�D��C�{uW/���=I+o����0`p�F�@ Tp�؏�c܄�0���2W�܌�����)�Y�2&�0 �!�Y_�B�
R�ડ��g������S��M�#;���+�VE]{�G�5�.�\�V?S�s�2D����>ǋT�\���-Û������3��\��iX����6:\$Оe�qК�(�����s�DW����ydKb0Ӎ��y��|�d��!�6��q/�&8e����7e���Hy�<�����7�����QAA�ܦ���	�V殛��΄�o���Ws��P�P* A��uh�=n����+�t��b�)%ND�cɳ���×��tY
i��H��1���}���?�ԥ����i�������=w#��o�Fnf��q1#qoG�/#��:d�|��h&]t����zl<f﯉�]J3��ۡn��X&��x�̷�'���P-M�?��9�/嗴,l��w��s��Ɗ�j�����f����G��ek)�E�5XJ����|(�T�xJ�'�����%6���U�����2��f���I���� >�26>���ۍ��9�nn���"�����K�s��ѫ6|�Oj���MS���Z�\��<A�����9aI�k��M~X�x'X���G
�1�A�T�LS�WZrʕא��/�����J�؞e��[������Y!7  Xa�}���F�>����22ǿo�QMN�o�Y0�����g���=UZꞯ_��ߥ�zk���D!�<YZ�`{���Av�bg���7N�H�Vg]��T�]�2{��ݷ��3�7a�cWȬ�~4߅�GO�!������R�c��I���3�����	�%?6�%�	^6<
POL��IO|�	��o��\�9K�j�J&�� 7v[o�A�j�Ÿ����Ӊ���r��{S`?����Z� �E�/R*º�5�f����Q8Ҏ��,xOv�C>49��>i	Mn|�H�����u��k�����Оܪ�9R`�_�Y�|��o��,��9@��*��wy}-^�N�;g�տ^��G�W�>����SȚ����wL���t	~�VS�_KDP���ADH�ټ�t6.!�8S֔ɘ���I�V�SD�<��U�P�$~��m��3��j��$i��݃����혞o��ٕL㙛wt��)� /���Q�-��ڽV}�54�2���mj	�EneK����cw:�ա7�Z��䜈�}·��Mv�N��.��"Ic���M�X������nߝ��)#߃?�+k�Ȝ���WA���������Ģ�4�@��\�߻�����|�}��P���_�Fb��DP�f�W�/� ��$���ƴ��'a��"���U�R!uIV�e�5��jf܈�9Px��`�kב��5-�_�9̵����.�`�����dx��&���rM�M��;E�L��x�j�C�ʐ0�ͯ@��9
>�ćD���&��<�}���}�m��3`��%�7t����ݚ�CPlۍ�����7)�X=�TfMŋf��8��H.�؅�(��h�8���^/�N���ۊ�ާ7��;�a-	��ⲡ�-j��w�/̙��H�|�A��!C6q�� ���|uox���:t��/{ṃ�>+*��^�LL���O��|<�� ���N*��W�KI.\_����K�e�d6y#�=(��#��퇢ɣ�q�V��nF��o�p�㯼��4i�엏����bʲG�Ԑ}�zy}k��z!��b}T�]��$�Ր��{FH��Y���4޾��
�ClrEӥ8_;�J�>K���d��ٻUNl;�� ���$�w_�c����ʜ��E(�殣w��(��
?l��c�?�s6Jp`���w,�����Q��y��z8�޵��7��l�=�YT��t��ĤΟK͌d����ј��l:��t#y���;kh �j[�t�@��!xZ��bB�_��i�2�`�C�w��f�����fW}͕�����ϋ����窝����ׯ�(��rp�d�ml��6����$�k��T��I�D}��q�$'�6��R���8���� ��.�:鰬�/�Y[!���&��.T���!v�O6^̿&%��Y����8
��K��an�jO�~n�	���/�1�E��|��VO>�չ����}���7�l�]H`�e�}�:5�>�7lUn����'4!Ⱥ6@D��?�jջ�f���x%>����^+�w��	#s|$;��sGs��ld�[������T� Z&�D�oƿ�ic�S�!<���@�q��)���2���� ���K]ގ㙚���#:�E�踔�P��K�G�"�>�O>��|[@B�Dv����GИ�U[Qr$�����;���/t�@�:��6yZ���m������2_$(�y���3�=��7��4�ݪ�l��mL�e�Cd+���ם'?}y̡��9�7��y)������X�σ���8 L�����g��|��Y���}��m9�Z�6c��+�`ҝ���k�Gʣ��RiR#�pB��H���Mz��X�o�#��I�r���afT��;����g},�@��<ac�� j�U���D0G�q2<dj���kϣJ,X�UT��Qt��7����S"T�"A�U(K���#Ó�C쉓'F��R�^A�`��6������,&=�gjh]Ėf[-��%�ѷyR�{��Ѳ��Z>�I�S�5[^PSG�*��Z����	�74s�E6UJJ.#�s�l|?�O��2�1~������3����e���0;�����y]T��1�NS���n붊#W����M�O�i���L1�&���ds�H�v`ފT��밼���\8: �b�+��/�8
F�;#Y��P�O.9Bn��e<.�_>ӈ3��l��ل(���Ը���~Ve^�)8UA�3S�9�[�VZ�.=s�j�G]�f\�?>�g�7��90��nC�@�ldڡ�eṼY4Z`�	�u�vGF,	`��8��V�@jJ�a3^�9Id��g/�71���F��N��x�*�&�]����o:pJ�dmvZ��w�?9E9�Ҭ.��<O�N����Fmߤ��G���	I"���bT���� �kJ��r�-��>�k��g����;;E��@�x�eq2����ߕ�}�ߟE�������޶uy��0}Pt,�oE��)�xsp���ʞd�T�p���1�Aq�P�\X�O����x4O�B��ϋw����|�m�rB���^�f{�mHm4��\X�J\�=%/Q��m�c�r[��3�=���\�^�°��!k�\~Z���՘)����7d�?�����a>V���2eMÂ�D;��B@V�d���fO��V�_ ���4 �LT<D�dK�U���\����2�ӹOK���T�=��̪i��L{���Kzc��J��,����i�?8�Q)��O�|�ܶ�-L�5���hr~����jZZV�4�ꢔ�=�j$�OmP&!H���{�쾴�}����m�;����)���C=����͝# {um��}�W�^��-��~7���_[������������Vۘ�����mw6�I�Ԥ}!K���������S
�U�X����c��Iݗ�v�3x�ƽ���(]�!R^�ߤx{X�:�H���p� ��&��� S�1m��l�6[�Ɔ,2�uG$O
�/�rٍ�8�Jlj��t���ن�ݢ9���)X�M	MT�pD.ғVt2T>����5����u�V�h*�����U��T[��=����N���ѢGF��	U������� }r\n"�������R²�'mxo"���E��kk��2�*�y	�2ָ����t��e��:-LbOuzcv~a�(�m��>�Z�o,L2t0N	�6�/�uu�^�����|S~f��2��n�$%��|	׹��S��(�9#���{jt\Q�� �Y-�q���"&�ft��s��3
����yݠ��r3�Cl��3���V>cKV>�磢�O^g�.V� ^�9 3��K��f���Ɔ�g��������e��A��x�%/*�]~�ч5.h���/D�G����b ���`s����q-Nu�.V�&��읋�ь���
�/��Ӕ������
ھ�Vك�p�NCqh�'3slaU��8�3.(�ql,X�����\ɵ��BM������d���1�tx��_wۑ O��q&����I�bB�P�,DV����0��,�ǉ�M���D @
j@��8h�gM��ua��f��y��Z�Ƅw�JU��c�t�W�6�L�9i�3X����h#]i(�F���1��A� >9SP�*1��k��ke�,�'x2�9:��7-J���K&p�g�t�A�vB�p�y[��6�y;Tu_������`���֔��b�X/'��9Q���A%l�|��m#�m�h��R.�9[����F�U���Rށ������Ie����'�!j*Þ܃Z����#�I�K�@PH%^��*hD�̝��wg��%��b=&0չ�y���S^t��,�F�oSr�2��A�^�����_��(�
F�}���Qe*S�c5�dd���,�"�O$�Mz]���JDX�
|-Dc�s+rŇ~���z����-�J�v���PA�5�I�/vHd	���!B�)Z�*tq�w��[��F3�y��B^g��}ָ�a�y'X���㛩�S��Y��>����~���C��F��r]�M�ȍ0�3��!��j�`�af���/K4Ѽ����CV�':j��pm6'�z2P R�>Xܶ��mʇV���+�9R�٠��)݊���f�4n��^��ih�M������vB*�@�$���]af�e�a��y�vڔ�>����@AQV��N�8�yM�hb�é`\e��(���P���8��K�t�BpC�0�H6�~2�ѡ���8:�r��PEiH�J,�_.�\�h��3�g.P�0y!�E/Cq����-4m���f��J�Uu�&�Z�g�K�em�׺m�@�E��hI��~t�U3��=?8׭ i}&V.4D��� kPcAp�2�����Ԡ��$g	�& ��}4"i��$��y��%N�X�w509����=����}��u��f�\xbsI����z��G?�i#ߖh��H�2S�^1vcC�oiK�L1�S9˓�E����'�ʒ��}ߎ��We����iS��jWۓ���@���@ᇩ)�m��ΏR�2M���q=4ͬb��ֹ���� X5y�D����Q�� ����~���%�o4I0��_�d��+�=�~��}ׯD/�6��e:�MJ��4��]��b��G�����<�#_�)�pJ����I�O�2�sP�M
�f��kd�+�5͋�#�pM.��U�1�fa��\~���K�u�f:xe�������;�=�\,�MM�?�Jp�ϥ�����R�q�,P禱P]P�@!0N�]�J�\Ə��-���s�v-Ӗ\w�J�սǧ����X{{��/
oeIVw�Seɫ���y��[�:+A�?��0Hֱ2w�K��&�{�o~�;�[�PEQ�����ۚU���U�h�#��V��&w��]��7b�C߮����z�bT��b��zX��1�3�^�=�\{W9׮\���#�,C�=�C@jo)�O&�n�`4�;�U�F
d������J����B�:���T�|l�"�cY����}1�c�Hb�#�9�{ї�?8Z���mz���P�g���Z��v!�t��aɏ�1��Q�d���'YG�f�����j�hW.��\(�3�Io?H>�ph��E����v%�����
r�:�=R[|'��=��!��н��-er���k[8�ϧ��Rچ��r���I������{Cd�*2��������2W���Ǆ�ļ����^I�[<�#bU�u�X��D`�G�?�)n��Jt
G1q��U?KS�o��|�|_3sT(�_6$هe��{��{EFWj�~��oO�1�����r��{$�&n���jo��I�7[g��ƙY]�ΐ^��j����g|{�yt�Ս�*%����Z�9�y=C!�F�or�:�7�8i��f������GY-�P	I���_�m�	�(xvM���=�B��4�P�f��i��	�|��>�����p׌�B
7��4�7��HӒn�+�,�Bs�ׯ�&���o)�`�����Y�Q�Gp�c´��V \��Mi0{��|��夻ߧ�t��>T��\B�������g__���&����+���)X%���Γr���&b!��8a����A(�a^�
p�	A�6�e�I��>�uOc�U�mr��C���ha�x Y%n�M�Uepp���9@�x��Sv��x�G�0}��Z�"������l�
ѽ���5]W�IFl�3D��ϐ*=���@�amrB�@/�%]^��}e����?��f��O�T[G������9�ɮ�������g���Nn1���(a��gd�F�"S]9���x��2���}�?��١��5��G)�P)iA�t�3��I�� �vS	Ҽ�8��َ']���9~a��V1����[������:�����ŁΖw�(Rdf�o�-��m�������
�Ηn��C$e	JA����x��J�|J����D�V쳊�pk��1K�u�4Hc;��I��p�N�f�t��^�3YB��_%a���	�H�F⇀��(|M���6k�I]-��S"����6�P�L8 �"e��E,�#/za�=Z�'_q�jѶL+�a:z[��ЈD�}�����3Jz��8,�����9����G��2��_��wz����}E'o��Ǎ-Q��ߖ<��v���+˕�Z)B�|(��+[=$��9��l�]ù�!�O�� Ca��DHEC���g����ӣ��ҍu�|���l�e
fx� �i���:�q
����@ϾW:�;��%�4�LEjQ��zP
�d&(��]�uy��.��4l�٢�6͂��a9�M�8�0Q}��v��j�������c��2�J�&{<䡞�p��̛�xo�Q������+}��(T<k���]B�k4~�����iZ����ʬ�.a�`�J�csOO.	�4Ǟ.%�3�QpU��K�_��y��v���$��<*Ǵ��]fҞ���J�c��d6��ē$N����V�Vj��eF-%f�LZ=�>S�>l̒��.�4�`��6E�7�u'�¿)�t:$����
ˣ�����j�'N����.N���zs���C�D�/��Psn40���E�aB����%~�ޥL|<�4>C'RY<�����t�c�=v�4���q�+}���Ixx������������P
*��果o�'��,ĕ.Z9��YS�K�&��k�R����{u��;�XΆ���R%i�{5�炍�_>�X�ʰ[�dM�ˍ{��J!�2*�E������6�5�K��)����[9�G
�h��4��/������c���u4�av���X��1��o�e�!���𔊮c�~��s�|��n�㭖V�u`U�8+N{rgGPW�D廢�8?�,��?��9�y�f�I4��Պ=Dk�n��Ȍh3��3��M�Ju~�`�e��=QN�ݒ�e�y ��,�͕_n�C0�NN2��[�S���#�v��-�y��$���U�� <}��?nRn�'�z�W(J��S!�Ο5�*W�'�T�5�an1��W�2E(]w�R B��~_nlym�^�t>W?��~1�uw[A����7��,BZe��� ]�z�
����<��
�v���1y{�<J�M�s�<� -��op�3��>}�@z�:�d�,�-�O��s���1I��l�A�*bEK]Ia�3���V4�OC
���$!|4�[F
g{[o$b�Ϭ��d�Gc�?���ѼD^��:g�K�]��9�]7aXńbOŶ��Ɲ�h�(�|���o	
7�P�$V5�ns�M���s޿'��ih�����n3�x�P�n/0*�#���VC3���!9C�&�)����j�yQ���ʕZ�F:#G���?xF��F�~�����W�|��*��xI���u1��|�Ē�0|�����H�7*�,��b����<�2���O����u%�x�J���o�Y6����:x<>�D3��2�s�5}7�~]��Փ�B��=�&�	Cc_O�N������NU�@
��;��{�¢k����O��I�9%G�Z���ͺ@D^�R1���#�R�l&��`3����B6 ��0�'��]I��EZ$!�ň�d$�s;�y>���iB��]���r�p�V�|h�f`���u�v�$��Šפ��\��"̵���J�t ���(D�N���6К��KAe7�߫���E�SG (����dfQ�Jr��K���+�QL�
�A���V� %��Cc�A5��r���{��萃��|�	}ؕ��{�DH��oi����Q����-X|�]ۅ@.�� 6W5������`���ʪA*���m��%���{D���>1�(���m���Nj�W��S�2�iak
hHmgE�h$Rڡ����[���3)"Ĳ���ka =�+�}�_[�D=�z���9�h�ڠ��f�_S{yӪyÜЬ� 2�@���2N����E}��M+��FF��Cu!�x�4�}8P���S��f��H=B��@����kRh�2=j�↷��G�Rt�Θ���F��JOߑ���e��@YF�u�g��jČ��i �{�@�'\���>���f�s�P.������A'������h>�м8��a̛J2W��v����3.���E1*��7n	�s���g�a6�D�<��NH���h<�R��s��BG�L�!��9�c�K�9$�XU�{�R���vw�}@�����
d��c)o�"��oS�s9	��*�AӉ*CX�yb��z��ByXI� r�8��Tza��� V@���"):����Ͻm׮��_�4?oo��[Xz�?_��O./,�|���f�-<��Q?�Y�nT��G8���|tt,8w%W4���{R��+#��̛ݑD!��C�7	�'@�6�#p�=��]~Gg(�`����|��K*qA/�{`�͘������?����??~f��a�����+x0�L��{_�3�
�m����s2�y�2���k?lX�4�  0�lla��<��=��x�	~���x�ɩ��L	�I�Xo��.f�g��ϻ?+����|e��a� �)��A;���M�iB=��V��ix��(���X؆���Z|�i�b0}!#��`�k0�D��T綃'U2o6��^�ư�d��q9w�9zlJ�����_�W�nm�O�������9����uY\ސͭ�4!��Kz-l�}��9H���s��;���<4��{.������s������ŕ#���C�.]biy��Z�~��j�t���ݞt�e�C)�.P#!|�TJ�UDH�)1�'Ib���fAb¦'�'��N@$��{5#A�{�EH㏇G�.Ă{���"�$��F�A(�7�a ��9>ʞp{F�kb��AX�ј����g��[l��c�K���fg?�����w��x`�X�ͽ�=��w��s����&�̠�_ڷRY�=F����b���-�~��[�/��=`g���G��<cB����CF*^S��� �5�NO%r��QɌ`�t�����ns�2Y<� sj@͂k%�}����̹J�85bY~
�nG��N9z�����J����)�ã����Srǹ�*||����b/���կ�;Ĩ��^������rS�dm����z�0ǘF����P-���=pǻv$�[gUv�<�3����\���p�����#/\{��������^W����B��5�w����rN�! ��e�p"׳|�f+�IA�-�g��{b쥓�x������
'��TG�*��ow�q����W�g�%f����O1�O�,К�I afh?��=�'�x ɒ��$�1�2L�K�gT��F��}�g�$.,�P3B�d{T�ǡi~�\K7�h8��:�=]��|v+�V�c#��� �3ɑ�����h9\g��X�?���'&'�N���^�>6I3M�D0�7;����H�
澟��2 |H�H�K�g�G�����=�� ��<�3}2�����EWN�8!'O���ׯK�R s�(��ݿo��uם21V��������������mo|�rG��i޼챜K+M�~}U�+Mi5����Ұ��,|�R�^��PD�C��>xϝ�ݳ'�r�p���c�M�W�p}��������<63{��k�gZ���V�>	�K�#�*qؽ�p!��(*8I�z}�� ����M< �{��R��9W'xW���Z7�}O�I��m�H@���$�h��L���_�~�5��	ϠZ��	�QZ�����˰�X�3$�Y �?�%`�Ӳ�F�g��Fr��<+>	���4X.6ɐw�g/��c�r�b	6Vz�{	�c�s��=����ϱn�y�����]_�88�,�331��6�A_��<�-?�~�ؗX���;]_X
B-r=_��:���X�2MP��|A2������ۃ9���(A�f;>}��Ő�0ݗ�eI���͞�>�R����qV�١f�g�
HL�{pr��;w���G���e��v]�������zsdrS�S
t�Id�ړ��%Y۪I��1�v��1I��3R.J	�����߻�S�O��Ё9�V���xނ��K��nw����3�/-=6;s�Ջ˫�ڍ�d���������XN�
[��4s���(h����N!����2�ў&!��Sk%lz�n%���6�Ām��$��K	���p=C��xn����c	ƃ���������|Դ�2Y�@�^��`�0Q�!��i3&3�ۤ͛}�%�,0���>PZ��i��%������NdV�_��5�7���B{ �I�äk+��q�T���7�����Ь,F-k^���� �Q��ܟ�,��@�9�y����~fN�:���v`�q��f��l�`p�@C3�������)�3=+Ϟ�̭�iA��(���>����g�X���9���m�0>1*�#e�ժ�i��ox�|��4���Y�7�=�v}E��kZp��� �$����Oi��	i���ؿ�>z����Y��M���
�Q�{ees�ʕ�g/]���ks��\�4OU��#�Zm�k�|��O�-�ǒ�8�|!x�*!�I��ά
X�"��NL�d��pQ�-�H��S0O�vJ@B��N���!y�<��^ %&Z�T�� O\`H�h�;�x)�Ic��'/1�DՃ��אY�iֻDmA�$E�!����7q��H�H��=KPf��a@>@�%�iT���az����{�h�Z/�sp��>y�BH_�S\~�����f�59���p��}��8s (��9�?��ͯ�g*�9�}ד�T�Y����e�a�����o��a�#�}�m�Y�1�:���9��|0}+Cq=�k���m��` s�9��=���ĩ��Ф5!��g�.-���L�4"���K}P>�c�##P\&9փG;$�(���oI�
S�Vm0ov�ɐ>�< �N�џ���s��3��r��U��y��|C�y��/��Ԧ�-.��:�����\ZYps�2�l��z��v7���$��ء*�������5���Be�+��zrH��8ۘ $R.TR!�:	LL0�`���kk;^�g�B�&�ҙW�ƀ�ω7s��m�(FTH$�^�D�%��c��~PeN�� NI�N~����1��B��6��Ϲ��h��0��0�Ϗ�.^K*Ӷ����W����C�^�g�3��`^�P����HB��?�0qγ�����	D4	�ty�9�	i�Zc�X<��y1p������y�=���~/���s5�Y`�q�6s$�c.��FN{ę{3���{��;��q��`�B�����>ۖ�(���{���CS	�"�S��L��^O�FGTr���#?��Q�2���*0 �zCdfvYV6�R�vT(����P sh�d�>>}���:7�?�r����M�����o80����f7��=�ؕW^5�����걍���V�H��L�hyܤkT�b
�nO���?�Oi��0�eLcP���H�x� ��ݥ�䶄
_�R�$�U�%|�Js�S"���]���E��$(�Ե�f�3n3&�$\��3-�w��q|��$�$� ߶�!p�8���c���'�P�}���0�=�F���o'���5�Ya���EV{�k ��3����P�co����M���}"�&���ǽ�=�/̝:}54j�4|�`����U�~?����Z'��ה��;����cu���s|��}yyU��a�S~��1�6�	Ӭl�S
�������ǡ{-��e�c0�ُ}������{�����(3L���v~h 
�(V(Ƚ���O����=���Y�T��i�Df����fMjՖ�ԍ��Csi{φ�뵫gO�����?���Y��8}S��� ����+׏^�r��/�rqq�%�Zk���N��=M��<
��TR�l�knpmڨp��I���!�77�62	C5��QH���Ԫ1!����ov���A�K��D�!��Ēj:e&�ݍN2L��zb��	�X�W�{�4���ה���T�w1�@�L���R^#�A݃9��8Qg� @� 
m���]mO2ۋ����s�|��L�az����H��uP��%��1Q��9f1� IA�?�4�W��̹/1&e<�]���{����
p�/�J#�[���t��ᷘ!�mx�=�Y���3��_�4�0,�����Ҋ,//�Ücߝ<yR�-��N'T��zG;\O�����\8�ܾKm����`��������� k���NZ����5nY�ʣj2��ܔÇ&�?�!�:<�	�����`��p4C���#ak���N�������z�\40_�`����oc�;����_�<���W���<�l����nw�P*K*�ل�����Ţ�K�n�B+H�;F���JEi7[(�k����}����]
��A.��J������/T�#A�N�bYZ�
E����P�X�����Y��y5>��� �p���(�D��@�<��'��X)*���O�>L9oT!3�=��<�g�/�=1�x�mq����8'��dmls?�YҢ�c� �9�3֝L�JFs�=�k��ٶ=��a`�>04��ݳ]˂���w���1���<�ׅs�6cF��&3�yr��
wY��k���c0G��@?�$[H��fx��S���3�C��1i�(�"��ҫ���M�� �J��͞00(���~.����nM9�<��V[��"��������[������I)g!��w`>�[���-Y��R5;���-��-DW�|����|�������������#�����ٹ�]�x�e��VY�h�6�G{��bՕb���v��O6{H_iī+#�Bi�l8 ��@߳"����0���Ä��~/i��,�"Ĭ�5G5�n���p0�~A	9����D�ĉ��C����W�-`D�dI�^��	��^ 
%d���K۪�۵K���x~��&GA\ )�E�����	 ����B�����a �߻t�8���x���8s��k�;>62wh�_�����qs�5�����H<'f��y��A��u% am�\�dahE�PF�e��r1���_K2����}>ׯa�O)�� �1�Lp�=X��H3%���s�{�+F0G��&^ o�9�s������އŃ9Ϣ������LC�I�!8��s��7?��Ȩ�����}�������}zzڜc��K?���U0���95��dhr �kiS���)�k5�V���Q�2I��w!G���C���C�K����������0v��g������/�3_����j��J�[��H�`��R���ȿ$  S��[��H\uãxϼ�������g�V�A|@Z
%<cB�ϔ�c�P��{�:f��!m̔rq����!d�#ъ%�����q�|�Ԣ/ա���
��	0���Za$��w�+��@ߑ,�n���h煴ȱz����m��9�f�2h�����VHOi�MJ�l�?�ҩ'�k�{�O=�"x{`��rofI�H=������Y\�0��'|���Z��<���I�8C�S���H���3��b����s�O�ɯA�������=�_���ǥD��.0S�A����H�o8��3_XX�:<Ãt��s��u�Y���F��zպ P3��Y(����a�I �,��H�8|�H�����c�s�%M{=٪T����u_z�)9�oL~�#�#��j7ճ_�ɜ�;����,�nJe6s
/gnc�^�#�vm����#����|�\5�+��t��3�g?�����O=��k��ݍz��n����p��@:����,!J'��0�Ԙ�y�<~�9��:OL<�z��D3���m�
D�Q�F�I�	�	��Hm�P�^Uֈ�t�-xM1�VUʒHܼ�אX4;�m*Zz�� � B i�����,�7��)�jE���&�Ѷ�Q�3`��_|�8j�4	���v}����3s���xb�W��W�s��n1�s�dNȤ��}J�Y@�y�Rt�������1S�9��S :�q]��D�e]�̑?KY��9�:3��>�)�������0�W
�~�����)���f3Q�C��`n����?�Ǉ�ù�5�|��Yu�E���<c���{�b�0�]���pc�^��о�3�� �O~�䱗� �'��	�BY �/-7̷6Z�Մ1�=� �Z(��j�Vz��>4��������3p[K������}��хK3o\�X�W*�J� �jA�2*H�R�iNlJ�B}l��S	;=J�B=�,5y���Ok��c�ć����c")�<y�p� �@��jK�{":�,p� �b��eO�:��DNU^W̌��f|,�	�ѫ�s@�ƃ9��� b�G� �CP�g�v��R��h�$�z*�R��|�3c�T|�⽒��%����*n�����'Kr��z�s�g�_3��r���7_��Q��=4��~���=���*>�'�b��@������|���x{��z!T�1��y�b���]���+�wG�MB�(��٤��{�����O�?������)��
�4�<�HF�ʜ�:�x��8O{��U�:Ƥ&�(���.絏JQ�Us/�/��eae#sK]m���k��ݭ����{O����];W�3pۂ92���?�������G���~MN�5{vyd\F���sԳh1�s�$Q%2�N���x��'6ׇ��	5�~e]����%/�� �KgJ9 p~\�Ԋ�W�^�|�*���;C�t����_O��g3�*�:�͗�����k�>�@�=�˕9	���b��Č��'�~m�G@{<���� J��#W �	��v�a$!f��1sT?W;�x�x�<4<���1 ?��=���n�\�=U����:2l�,����� ����2	��0�i���a�zV�?@X~��)�,[�����Ѡd��Q;��O�{�"��m�`^�|w�����U�̬0�ܡ-2������c��,�^ő�LF ��d_��|s��-�W�9��ig{��	��<���.YYYт,�b ��;����ͯ�b+����#��ԑ��u��hHO͗s� �PaHV�~[ڝz�γ'�<}r����v���m�_������'W7�F,��+=ׇ�ۈ�r���[�w��3��a`�F� 艥'��Ƅ���yu[,P����4��ų�BOoK�Ԕ ���OP����Q��.ڜ�8tO�H�Ʉ�w�6	�:�E��g(��C� �7���Ǌ#	x�>ں�^�	5��k�Ǉ>@�"b��I����#! ���:6YD:�:/�e1d1H�y�yjvߎ_�H��nRY`��O�U��R`>� �γ�kocD Y�uccC�IR�6Y�#̳ ��\�<sb���U��k�m�Y��f��O���9���R�&���ԔF��z�r��ȸ�^jQ�7����y�s��:��ZT�{?��!`���G�%9s�J���h�hcj�e��Z]mk��EV�����]��oz����ߖF�`�ܒ��M�np�3�����Am������#?q���_��rV�u�u�3pۂ��������ٕ��o#���N܎h�@    IDATt���J،�$ą�U�RB8\�~3�c�����9%AV"�9		��U� ���x"Op��$�.QuIg.���������@�c�v�'�vA�E�=�W�R��1���9�!�ǫm)u+��
VJ�$�&�`�E&�`�)�S�4Oo�����a����y�ƀ�O�4��3E���z0z��p��z ���a�d�0���lyS� w�?��ä��h`�6}_���C3�{�׃�6��{�����[�47~\*4�tR����{f�k2�;�`>77'���ѭ# s�~�ذy2rj����h�a�yC�R�jE�f�9e0���qjv�W:�_^*�P0�[�TM�8|dJ��67*r��UY������1��|GZ�%��Վ�/���ZM��m���}H���ُ9����}��s�iO.�-�|iii��?��_��_<��F'���bOˍ��Es�V��ZIU2�1s��wOHcb�E���ܫ��̘	������hjr� x��6h�z��{�$0yG3��E�%(��*U;�H�S4.?��]�5������q@<���v�ԱT�\�" {Bǹ!���H��?�c�,3�q�A����~r�<�C�À|غ����L�
��n�����"�����a�$��B���\��5�
>�J]�x?�sB��t`�����{�:�Y���co|f�9��_����;�D�-m���V�Ӳ���Ql��Z9�9$s���t���Z ��>�]2t��7��9^}0�}��Ό�5:>��s��Š~�a������ΎMLh�+[5�p�T�5����o�O~�'?��^��
t�ЬotenqC�Iۣ���4����!�)�&��/S�M�ؑ\���nznK0�|�:���럾|e�U�~I�T�B)/�т��N)]uQ�w�	!4,^�؞�yu�?��`��qV�٫��{c����}��<&b�"�e�6���Dr^z�j}H�֫��]�53��׫\	f����ǹ'��a���_�j�'|�ʱQ�%`���W4�G����~��<�
�r�����d&h��3� p=����XM35~�������#ٗt�$F��W�����{�K�~��@f#�s|+�}M3����ǃ�������ݫ�	X��� 	0��Ű4\�P88My����$ȏ����b*�>��g|��5�p��x���i��z��EM�8H��}�U�vi���܂���qا�B+��A��9��@¬	*9��A��i��)�y�0!�
�����P�Fۉ�[(��	�7>��}�_�~]y���?��2�)�BxZ��#qL�*27�.�kUM灱�^��|�;B�����KgN��}�rk7�b;����K_Z<������\��xa�c��FF�2R��:�s�`�"�>�1�j�X��%�ĆD"&�7�38�0���,4.�X� Aa�*da���t�)���w%��k�Tݔ�}IJU���Ơ5 HIdh��gz������ EU�ys����ZGp��m�h��*]������5l׮��&�V��� -�E�>׃�$P�sLX��W|GM����7#�������I����?�Ü2s��d� Ks�3��!����ד^�^�iPa-1�x&�k���s����g��=����ُ�32l�k.���ٍM}?<���4;C)��5!��v�j�j��fI[[_O�"@M���٨V�͜��{
��bh�ߣ�7J.Ce���o4'��ă��3c�zM��׾��rϽw鞹v�2#p:V��վ̟z�)��V�w��=�?�9}b��I.�[�K^:(��Օ啪ln5�RE��1M(��W�h��bN��/�ۻΝ~��ݹ���n�>ݖ`��y�_��������]�ވ@|��9�XdC�>�>�C�b)(�ϒ<0#01�ǜ/�����U�9&P���M=蘊`�&(�{�=���I�TR-Z�4�g	�y������
����2�e�Ux���?��'�ҋ��p�`��ML@i����L����6��%�A�����|#�6~��K5��m��1�����}���Ҩ���^�Ǫ^�l��	bԆ[�*QƼ�/@�닶hn�\�	 �ӟ���L�E;�_:y�;D3 䱶��OL���"��m����x.cov�}rn����7�	��s���7;�FÜ@�XG�&�S�No��$ �M��v���'�r@��W������ȋ^�"y��Us ��W��A���L(�J]._�,�bI�%�}�"����s�)M.hQ_��!�olvei�"�u������ `��/�B�Ljy|��S��s����㹙�8oǾݖ`�G��e������j�t77"�RYJ弔FP2<R�[�1<Ï��D�	���)|HL�����?0$YC�����ܴo'�-Gޘt�^��1K��R	a7j������F��>��KG5� �U1�<��=@69��s�H��9��%p=����2-Gn�39?j��P���'��k��3T�c�L�W�z"��v`H�c�������e��o̳��o��3��U�_H�^�5�"��ƍB!��u�Za��ŏ�fp=���x\���� �Y���s�t�w�^�����2?�,F+a�Ԅcq�m��!-��@�F��k���F	�7%s2����i s�h!���x�c�d������t��-���w�&aNh'�P�1��r�wȣ/}�����n_�җ�F��!dmyiUMȼY�wd�ԑO���:�R|)�
�"6󎬬�̷*H��� {���M3G�B�+�����챷:4�����s�nK0���������?����^~TJH�2
�M��yN
�;!�Z��#0�A������'�Y��/��'
Y 9�Q=n^��I�b��g
�f�fk���㐀��*��(��h����xɓ�������^�C?�t��\Zm#�͚U�B�(1RR��d@8�����(б�C�`�ES=�M��%�Oس �k%<Ϛ?O��a۱��\`�u�?bI��2T ���y��B��B�,��`���vt2  s��������!��D��S&m�ϸ�E`���������ۢI�k^�$�h�,k�����\�<�zߌ�1'�w�����Z�m �K��
?����ψ��}����дx~�ͮ{�/zv�]w� �P���n$j�R�,33�4!����wd�ؕ�����7��B*�]�)]��Jr��Փ���ln4̻�`&�(�%��:�/t�\����c��M�����c�nK0�����w����qm�y ���h9s8e#ې�yO��G�Ul�_O�<���ޗ���艩�oX{	�R�'�ۙ���Yϊ��m}�g�9���j8��zMǵ����M�U��{ �%��<x��R:�s�!iMu��a6!Y�}���
�A���*Q�L��d�w�%��Ԉ�`A	u��~~��\G��e�1�;�&a6���dHa#����G���l�7�s��G'�5'd����{���aqƐ+��ܷE���Xg��i�A?���(k|Èfr��T�~��sGI��Ҙ�4\ֹ	��	��:�h2��VOm����;06P���f�2���%s/��?1�ǌ5{���9��/�iQ.?7x߬���ٳr��wk��H�(O?��4ꦡ�d{��+3����q�ْ�=�׽(�^����N_dk�-k�M��l��&hP(���*�w��̦�mJ�ؓR�7{��ԻOٽ���9������������?߬vvInTF�Fe�y����.�z�]$`�RW��5�L���	�Y�Fb��_�u�>�{cа����xL���=@��۸�ȈU����S��&AMTttP�$�?�>�cM!�v�U� lh_��;ih%<�}_�l����<���E�0 1!2:��� q4B�f�d�23�*��a{�T�������3k�{�`�n�y�xr�:�����k!U�>� �&�� ��Z�/�.��M<��5��<�H����Y�ϫ��y���f�ϡ���d?�eb|��`���ښ2-�;0EH骧�gsB�%5&�~�\�9HU����'s��%B�0'�|߾��裏�9:2}X��VW��i�����fEU��N_���2V�K��"�|��mo}�&�Ԫҽ��%iv�R��e}�%[�Y�@� |����\5��K}����G�x��S?{�X������~���������?��5�ԗ������9dzc�sj�ͻ���̵9�� ����fOm��D���XM�x^��sӝ���0��.%���<�XX�K���7���$7�Z�##���A�$�4Ýٶ��s|{��솶}~罼c���	'M�C_�$ �0N�p9���]�G�*J�3\���}��~݋A�ϙ�/~/��SSs��/l�?�����V^z�����Z�s�5��:!\(�X	��S܋� �L40����{��vwF0b�9��\�����b@�jPg��k~�dn{֞�ϧ�E�f!����4�̗���1G �cǎ��f��4ip?R2�3|:ט>��f��"'�����`[���-����׼��)�k����c�
e]���*�瑗"��My�_#���o�]Ӻv�-A�Y�ޒf�/��T����^�v�$s ?�^U�t�us�������L�˯��?�ڸ�����[?�G�?�� ngD��22
�RO��$sK��C^� �gmv�� �i��6�lG8��p�,�;$�	|�li�!~yb�c��6&s3C2�$���F�������z���z�:P�҃~�/��wHZAI�0�m�$���iצ䋿��h�'q��Him�K���Aߠ�ĵp�ٳg�JFh��E�j�?�x���6L0�6����m���El��5�?�9�;�+o��5�	ڠ��qjJp-���W��w>�:搹סY!s��X�2�i�s3(���V@>�!�bS��iu
�����@)�S�s�qp�y�gP��?����$/���c�'_[ {����ʃ�J0C���zLa3��'��&0�.y��_/�fC�M+���J���:�9�{ʄ�#���yL>����{B/ �(ǺQ�K����-٪4eu�"���:�̱?ZͪQ�]���?{�]���NJ�[cEn;0_\����g~��?�����ے˗L2���E�tu3��*�������%%N �C���+&[��b�N������>gq�ޛE�����AqL� ) �EL"�T6�up���Kn^�5bcĀ@�{�,��qB�{l��P��U�q� ����sC80�_���6 U��
�E�h��z�ۘ�/�6LR�d���A��Q?�����c���c�ׁک�ir������=�j��Jz�g� ��3y��x\�3�W'Lg"!Ȱ/H��U�~�����Z�<��=��A	�<��g����O�1W9����ve���h�P� 6s�)���	٣6��M�F��׻�;�8C��q����{}�9��o��3?g��h��	��6�yF}`����/}�C���n�PD�����"�m�5�Ri6ec�*�F[J�S�J�����\i$/�~���Ջ_p�#�\�rkp���������������_|���4`{�d>�8L	��I�qh�?�$��z�+���v�˺��z��@��D�>�3<|�|�\\R������I�d>�rI�j ?<�)=ch�\!ޔ��Lޣ]�9!R
�2�MusC�c�1G�@&��G�f�B3:j��$0h�aB;C���PC�&�ٞ���J[�C���G$�k�=���y���K�6g��=�*��j�~������v�9�D0�s���x޸/8?1s�q�s晃nK$��~�s]=�q|�~.��bZQW�-f <��ג!k�����s��aN� s�?J�wC�T�я���ΔX��K�y��1��D�8�d�1OP������/��1Rg�*��#��HE5��C>��{��^h�z�T���K����Z[*����m*���F$�1SZ7/҅@��RN��4"�����o۳'�����[�m����ß�����矽�w�͎�f^6I�6��܃�˫�<QT�}H�Wnf\O,}Y������#�𿳏$8$�S��b|?<A�3����9t�}Ճ�;�E��qມV��:�j<g�Uγ�1�ot�cw�����n�t�=�� �y�@D�-�O���ߐ|��	Ц�;	:�q����z�Y���ڏ�}��2?_~�y�u�3���������F2�d����9�%��7�q#�i��}���yf<������b~��$���O��3= s?�؇a�����G�ǳ������3��|�!���!�9��r#��U���4��j��v.�t��L0������;R3��M�@��A��^j^��B8�˕�5=Cc�L*�Tj�fg�@<Υ�?�O��~�=r��-Bӥ;Gꍾ4��}�-[����oJ�ޒr�l���2EW��H��:�Iq��g��������=������ڵډ��S������сgT%�҈9*Q2�������o|<�y���0B����=X����g,��|Y Bb㟙�UY�"~���M�H��z�TI�;�	��̇!���{�u$�z�	bI�*C�éR��O7�H���J�՜|	��$<����F�9�%J��Q v�0��m��$��\�D҃��e ��_J�\c�n�������5f&R�a,Ge�+�#��7��	�Ms�g�	�|f̜�n�K/uf�U��T����d �	����Ls|�؎����b�������2��i�PLeI%\�]3�����`fw|����t�7�*/l��	Q<���%Β_{\�q�/u�����D�g=���j���lT�t~�4�}(���
y��W0���i)�{�ˣ7EAE�ZKdm�.�fS67kҨ4��+i*n��C��#&��`�/��>s��[�N���\��/����6/�^]��S��7��ry�ͮ�Hi,s��`KJ��z�1�{���[*+O(�yJ����&�mg��I�cU��b0�ױ����0�L� dq�f��m���±VK3HE��D� 	PEO����k���_<D IHR���`�j������(��5;��g� ���4�yD{x���5�|~s�qs=�� c�s���1��K�À�{�{ȃ�q�F��K�25*��X�%��^Hl�C&�����^e	�W΃��a6m~:!��$fT�f���Ï�3;������s|�s���'I���=�7����-C!�݊��w�$�s/��ttK�km�S�����]��j3�W�r0	�޽������dIu��F�K��	����ʲwOQ>��>tBJU�y�z�+�VN�+uiwav���</E)@Վ�`^*BK�h%�Iu��<u�;OL��vç۹?��d���,��˟�����.�_��5�6n�l���yn:&�2�x��I�I <��9_J�^�o�c�����F��]�Ս ��� ��Y�$�i�#@��̑��Tzq�x����jD��5�=��\�Am���;����y���Z�����*�a�ޣ�ƃ��01],	 ��\�d 10{���G<s��^��Tc��^  z ����/���%G�5 ��K���gT!ty���=@��gp-BӼf�}���42��� �6s��pl�'�ܟ!�r��M!6{!�ܛ�<#��� >^�d�c0���v��zHY�ܘVs���d���0���=�L���̳��1.���/-�2�/ 8�)g���!�:K
�&I�D�e�DA�����SJ��}i7{�j����\���j+ˠ'���$ �<LA�@!m�������G���齿u;���ַ�����������>=7�rg/_R����x�f'��{vȕ+��Y4�#�փ�'�<�0�����o���A!�{⤑Q�\�܈��s/푨K��    IDAT��d�L������d[��0b�iT��؂@�t�$ޜ�/���z�#H�v~��a<� �3���A8	D�ǗY�C�b�o���W1���g���3�_}eI��?{�$�u�	��>+����аC�)�^t�fő(��Hifw��������V����@� ,����4�Twuw����J�߹��<u�U��?*�S�޻���|�����-���H�����w�y/�d�����h��5��j_��>���U�s�	$!x�-H۶��,ڽ�t����ד���(s/�:�̫պ�qjvM�S,*�f�����}I~y�6�eG{ػ�<�f�?]K�c'_�g�<a���8;��e�XJ-<ٵHN��(�V�6!�K�Z��lL���Oʥ�씶�H&Hi�*�*��5��/h��b�*S�Ҩ'$K���V˂L{u�ؑ�^����i[���� s%�gŁ�S/��߿�;'�O�ođ�-�`ovl^�ٕ(��L�,��	$�%����5��ؗ�Z��DGA7��6x�s{�%���K�5=��=���	^��-�7�"��K,I���0w4U�|&Uw��jw�t5���l��g�3c��>$�l��ēk��g���vt&A�}v��kJ8.��q_��s������e�,��~��v_�>�~r��Υ���VZ�����τ3։�2��Y�$n5>��v��g��N�ؗ0Ϟ��g,3���-ݳ&,����3����{���g���� ��:k�\]rh�\9�S����d�u\�p���I/B�f?jahm����s�!����c[xE�uh������ᴗmS D@���l�v���N�"�L _��G�ҋvJW[\R	����E�񩹂�I)Wj.�;�챶&�!�C2O��5/t�������Jϕַ�=��w�y��;=5?�L�M�TS2G��<�M%KH����O��F&(D�˃O����4ɸf`��i+yX���e�=�I�L�%��~K��h�`���K�O����tq�'�j|"o��Dh��L�;ߖВ�//����9wT1Z����g8��Vb�����n'�j�}	ѭ����9�}�d�l<{�art:�g?#��pc��6J�dZ�e|�*yv/�y�=C��k��ڬd��� �~I�I~V�OM�a�3  ��K#�[&�5�
�]�d��0\��Aʠ��b�v7��g�,S��H�d�"���e&a�!�c��h3��p�B�P �^1����%��f��s�BK����5B8�������ң�̕i�A���Q%��c�����g��	��Ro������q�&ٴv@h�����,�j23;'��Y,�ejjF��d�t�	+XhH4�Vt��j���;�:����+�?+��}�O���yf��Y�%̡ʅ7;�&���_6��JX������Ԃ�=��fq	/%*ז�� �~��J�c&�����0�חH����M�t~�y�m�g����]Fͫ%�H:BP�\s�h/'06�̷�Dx]�:�gd���ϝό���L�r��3W��/�#�ӳ���g����WJ��C�QMI�_C{��0_�l��.�Y3 �P�%6J��`�&�1�U��%���ު�	��?�T�l���������f���l����L�����iJ#;���_��s�jv�s��Xc[�#���i��"�)A�j�����zę�Zp=�$0\��_�wN����a� �C�βŚ�!J�H�%i�?F%K�q:ِ�>r�\���ȱ����g\b���@ �1���Y�UQ��%�qu�k
�E\�Y���Խ����'8�R�s��kŁ��w?��?����S �l&�`�Nb90�����mr[�DؗJ9����J ���D��Z�z+�X�� �?6�� �J���m j���yKM�d<~���T���bf�u�
X���hϪ)	�/Qٵ�������5�����{�_��q�@�{� �sB�����쪮4,M��0)�s~GOi�������?>��i)%[
�6����:�4����&�Ai�2q�P�gnt�OgH#�@��y���	ˀ���\�0�>�/�(���U�x��g��=.q��XOęc� r��E����M��,dʪ5��RȾ�~�&����瓡iP�G�<�BhҸ�lV#@�W��ph����Mm��M!�nQλ�t����e��5�k�Eff*R-Wt�鬓�gg�R*�T3���u�Y�K}5��U�n�Hg��AD�H������F���G���_<����Ε%�Z�]3�I�_�sn~,�U���#���D<�����4�b���E�O.aj�Q�HXF�V�WQ �vOܪ�z� �^���X��g ��9�S����(�4�NP�N0�x�'�_�ti�5j�,HXI���ϱkd�;a��D����ao��P�y�	JL��>��%�O��io�=�	��rt�xQ��x<�O�+��(��yV-op�0vD���W�����\eיaR���\���>�d��.���^@F�����/G����
|Oov>�0���d�W���L(��d��wv�t�� �]p9,�R�<L�ڜ�P�~���������\z�
���K���	�
��:r���5���K/�%�]~���qI��R-�?`�T�%YX��x��c��^����9�Y��!Ǝ��������Ϥ�/e��� 1SKH!Y�Te��"J�w�w;wE���h����ǧ�{����� s'QփV�
��}���9���������j6�o%�( �����6���'�ˁ���i�����zJ�$>��톅f��`,��^�z�85�҂9��ϨqPz�z��X�GF�g,���-7�d}����(j	4��Jf �
����@ZB{֗�ҭ[�֔��̍ݯQ�
��	#�}�{�ڟc slǄ��v<M�	`i��ѐ�h�%@��ҩ� Hw��k�0h�E]��Ç>�;�D�g�m��=���6��??�n9&��Z�9I��2������2Z�ܙ]�fBx���`N��$����0�-��g�}gnvJ�F�6\�L���+���_����<�c ��|��m�6����s�;S��}�V�����t^�媬_�V(��d��A]���4� s��jv֕wg���]���$�I,$�B"��ǂ�z�2_�5�Ej3��N�b�7�xb$�hLAc��NN�f�X a���ߊ��F�������ޏ�jg��P��A��O�檚})����S�u4ir�	RXt \��l�'�� `A�ﱡ�k�v��,��<�`5~�� �YF�;K��[ܒ�����%�:���o�9~�K|v�VL@���,��#a��*�}��v�D1M����ڳ��ܐ`�͎�rf`cB����8\0F;��_#���T�a�c���E[��,���82}�q� ��8�-��3Aï�9�R��x "��������q`�`��^��ޟ�%���,SGP�>�y�co�yK-�1:�s'C5;�-�5H�2�%�P,j� ��jH�B��&CӚv�0�;��{�cq�aة�gq���wH�n~D��׮]�dp`XFFF�}{�I&[�mHG�U1A}������k5��b�"�DN�~�����\Zҩ@�o�,���hxZ�`,� �=��c\�z5)��y��p�����,A���F�Qh4j�F�V�'�H2��awG��;:���%8_Q`~p���߽��{�8x��bCH$�9�� s8��V����<U��Q��k~��4%c��ިg��f ��( �}�&��(��7'L���$�L(�L۷}��Y�DU����7�cF��ǵ�-o�#|�u4���z����u�sh	\ԘI`|���q<��T�.>�1�6�ϴ%�p����0�Z�����sD�K��J��!�϶�
���'=��   1����\�PqIc�S��2$QJ��MӘ��9t�c*_��	�(�L6�X�c������}��?x�Mp�l�4G��$�/�B���������8	l�3��~�[�N�Q��r���ODm�W:�62U� �~�+�bL/�� �k�BJo%}wf\x�����fhhXc��\A#&�ᜀY�$S��ѭ�������?+������sP�;.��y�\[B�9s��K�
�RC�:g.r��Q2������H{G�:�Af �>C�ޤ>ժ�~��4jiH�hG6�CC������_Q`~�Dq�~뇷�?px����m�)����lG�X{$�C�ĺ+{��(i+�����o�A���8 N�p`n��p�o���R�0��?�!!��V2$P`خ%F��o%�c��e$s�ς	>	^as#��ݘ��qȶ���7�G;���y�z���y��Gb���ᳬ}�2TL|F��TS�e�T�P@ ���{��e2��=4.�^Wp���ߣچ8f���g	Y�C{w��kc(���o�������U 7��!��L���뵚^[�2&4�`�0/49@};��w���5�~=�V,S:����{��{� g��c����|l޼Y�\����U��`N�[�G�P��J� gϊ�y�*�L'��d2���s��*<�Sqٺu�|�c�/��C��D�Jfd~qA��g�I���:s��Ieeߛ{���q��g?-�¼�w�J����^�fP�i����.�R��y=.�Z�|-�\iT�a�E__�tu���a�=�ᐚ�N$��G=���<�&��}ݝ����&8���YQ`������r�##�;�U��&$��J*�Z��s๴`��6I�@���L�O��ae�Hˈ����U�x��Ml�>�U%[�Q4�-�L�1m�Qג��y"��g4��
g�����U���������7�c56��I���hz��^�(�!1��[��؟7˰X g[>sE�<�U 0��m�>Ӷm�@@��pPI��E�Yb�d��Ľ�)5e�f��Ip�g2Rx�]��t,m�l��=�<�9�3l�8'h �}0s��@b��9{q%T睊 ��IB2f��G2鴶���C� ����yX05d� �}������n���#�ǸN@��b�x.��c��t,4/`��:���q�Qދ5<�>:�e'Ż�H2b^��%�E*�v hJ��'�H���"��ԇe���嗿xB�}�E	���RmR�"U���׽� �ʴi��ʍ7^�ڐt�M*�@���%�
$�,�UW^$���椴�Pf�V�ψk��0ņ�IooNuК���?�%pN�hbq��`��RZ̿�����ގ���rooE��+�N����u�����z-.�dB�0�ɘ� p�=�a���k:A���*T6���Z;H< l ���an١l쁷 �o,��L(y�̆��'J
��q,�z�Nm�Jz;.���e�,�[��WA+�	5,�y��O��)��({��|�=�1D1���[&��c��ߟ�-�g� p � 'ր@`!��=�@�_h�ը6�[���X,̤�ғa�2��Czĳ �̜5�W)9"��7|�L����%3a�4�� �h3�H6���^c���Ը0�w��1'tL�R��K��Ji�̕O' �v=�~�̸�Q�-��cųG��*FF	c�Ӥc�/��>H�h���x}w=T��eJ�^�D��q��}��Q�.��Y�ħo���r��?��}FR)�R"WV?%�;5��5MH�@���9zL���+7��Aٰq�J�'�O�\~A���@�-�6�nx�$���N�Hq*vD(aOhɴ%`�yo_���ձ�
�h0��UE�t8�K��xyM�-�����=���J��kYQ`��#���o��,��$�)u��g#��h!?rђ�=	�%���u���7��wT�B5�������#����T�(�}��������[�'���( �ۍ�l�Φv�pv||�
����;���ܲk�$�F=���6|�5^fK�O�\�+J#���9���   �� G{�~�.h��l� ds��v���� N��%Y�"�S�C
F&�x�k`�G�����-�7���Ү �
jV��~���� �O?�?����1.��a��Y�c ��e�u?�f2���Sx�׺�w�\di߫3[�"GG�7k�s� �`HT=^m�P���+5G������ �N��*��4@m�'�^� �fCj����W���1���'���=,�F�Ŕ�BXR0W�N�H��ߧ�iO����/�$�}�{墋.T'����ezf^�2==.�DIn��*�eb�f/�cR�_���M�V+�s���ҷ�H��b���2��B3I8J`P��:2���>��ж߆kV�?���k~���=69�Z'�d2)A�M��uy�B�t(�c�Y��'�$^Q �����j#� ��s�Rj'�3 >�,'�EI���3!>�X��g&,pr<�¿�Γ3;�Vb��lߚ`:G�~F2H�V����|�����9X�9�ėV8N�|5Wd��_ۇ(�?j���d4�0A�u$s��.L�ki:H#�Cʦj����$��O P�&�3�+j\�.w5�Ѧ>'��0<<��Q�c��¼�}�X���*8���&���!���y�c���� �/`�0w����1��&bR�ja���{�݋���N��+�V�٪U91֪��u̛c��2���Fz�s� �V#��9����l�̼K��!�N�@�TVɼ�++\t�|ዟ�g�]~��{df��$\!�m,�c{z����yy��W��/�w��
e�ff�r������ѣR����.�ޮ�L�MJ�G���Ξ(��訋�q���m)ٰnU�)���n��E���U���xL��Z)��e�������T^[Q`~�C/�{��g��s�= �ݞ=��g���Q\Wsӛ���x�i�%l���8J4,w�p�}̀Ol��1%Q���޿��Q���3 �m�m;'7k;�g8���N��kH��s_�a����oC��!1�Z�����8>J�'���p=�'0��tI'/���V �B}���kH)������`�H0�������x��P�%��=��j���~�4*$i .4	x���1��6ू�ڛ��*���|�ą�\�Ҵ������d0���\���ﭩǩ�V��t����Һe4����1>��YU�[.�g��̌^_w�9�ĩFG	�t��lJ�����C��?Mk��땪�^3��>��ߗg�{Un���27��n�ԑ�LZ�#�@8����!C���){s�r�;�]W]���<|T�s%���Z}A.��Y=�#c�Ƥ��'�&G�I�8������ڰn����	�
U��s�c�0���J%n���_�K �[�������<��?����-?_�5�I�T�$�\�BN̗̭A�n����D��ԔZ,#����yUV�s��� lJ�O;j'�ˁ9	���\\���aX�yb{�,c?���`����XB�gR�n����m�T� ���#��b��Q�a��֫�D�_'����
�@�%���N��)�N�� j ���%s{U��5�er_p\�����v��f�$+�[�X�&V���S@�{���042:?Ʉ�B���T�� ���.;��a�>�&'���a/7& �
����y��=4~V[e�(�\�3ϗ����v���9��=Ƶc�]?��P2��`���H3m�xU8�U@h"
���qK�ܹ�-��3e�RE��䪫/�������;���ĤC2�6�6�
���١Q��l��֪F��[d���r���J[�3�>rTf��X.I�\�Ӷo�����D�Ή4B�����_�i�zI$��.�dR��U��?��RjO���`�r��qg_��A��G���>r�C�<����@�<p��TK2����1a��:d�)I`|`����q�xx���@BΐD�0�����^����b�+�T� �dc�h�i	���N �o>�Y���=���2Q��{I,��>��kd�/     IDAT|i�W1�/Q��[iܪD�Y�g��]�l�glh��{�F��9�`� ��6m� ��g�mȐbx.Ӯ��Դ�S2��ӽF 6��8� Ζ�Bl������x&���Xq2EtLc9����^'���츆	J�x6��x��&����aB8�_���ٳ�/��Q���w��oy,��L>�v���RѾ�0�.`�^J�����*]dt�ﺆ�s���1��2G�<kU�\{J�~�e��Oy�1��O�U0G�S�����s�I{GVV�q&���Ⱥ�����aioG8q\��OIai��2;=!]��6;>����1�����B�i�l7�Q0w�2bМO*�+��N�����Y$�K�Q9�ם����ьȄ��?��m��W�d�h4R������G���b%&� �}���#�k�wÁ�����W��;	怄�7jJh�!N8@8�hǅ�8�ڰ9����)Jߖ �_Q��Ql� �@k�L�Ǫ�ض�]΋/��c�D�2VJi��1B�8��X�c��UY��ڎ'j����ϳ�f�����<Z��=�m����w;c�5��O��H��q=��;ڧ���9��!Y�w���x65\���m��1�`��˚�6�5�F���9a*PJԸ�#�$Wf�C<6�%���Χ�?N����d��m�`���kA0�������Y�+�bMH4{X��7;5�;0�˶m۔V`��Ų6O� �4����0λVs^�ʠi���"�f9ps���z�?A�F\���+Ε���zy��7��?�[��5���s`8�ԹK�⩹���)=|���t<_�ܧ���K���2==/�yik�ɩ1I�����&���I��<���%�����I$�Y��k�4��ktvv�dq�K�S���|��%C�b�� �Fc"��^��C�z��h4A��h<�����j&��<ޡV���7:������k���b	��N��ov:��P�@3��nn����An����L{��
�B��]�Y"�t� $�m��|3|��\8+�(����C�>
��(T�\- ��[��mZ��-���,�e5�����>�kl���g��y�,�rMm(���ҥ��f��(������@�Q�f����g:�kv�жJ���:�mذA�cϠL��P²�D�m��F�˸n�|���$szL�? V8��V�
���{�9V�V��y��|x�CJ���{�&(=K9�9��g*���2���oJ��}���=��H��}�y��c\O$!��X�Gy>zg[���6��d�&�&�ɩM���� ���3P���Y�8����:&��c"�S�/�"]a����ҭ:z�߸��{*H"��\p�Yr�{�-o�uP~���J���lHT֣��ߝ&�f�I��Ωic�K�T���|\֮P��릦甎��ĚlݼQ�=.�ź�*�FT�TA��svL��
ƎV�d��[�{�(�&(
���` 4�0=u�u�k`���iT�.*� ��(S[*Wk��L*�ܳzͪ��=#����0?27�w�7����{�TF�xE|9�-�[5��p�-��=	1��*ld��UJ	��;�6*6�=��a�jv�|~V��<�ش��a���r�>X�`��L��Vb����6����h+}��9��|>`5	gD�>K��dK`��������m�����rL�`m�|�3�oQ�a%�;5E � %�:%8��E���\h�e����_���\��2뚟�*L;(�B�I��O��U�V�wx.����	8s�������"��}�1k,u��s�ԑ�k0�5�3zF_5�>L=JfgvnN�OFm�4a�̗04�Τc�Aߞ��~2�
e<k|�B�`�5��9��C�L����['��L�ǌyijL	h��t��V��yo2��d��t&&[������drjN�����4L,�k(S�9r��9b���y�Ž�J$��I6mY%�@x������ӫL#�n�,��s2;=/�JM%k��2"����yѐ��Ns8�1W(tM0<��Ӄ����8���}���)�$
9����=ǾJ�T]54|W*Q�Zggz���J�mŀ����U߾�����*�@�ɴ����s�4m�̛4p>���H�v\��р�B@��])B\KBI�k�T��py���&Ħ׍{��A��,�J'>�'�����|��/�,�d�ن}����۰�����@�>{-��}�%�Tc�Z���S��23��u�eR�7�7׈jUz��k8&���N��W8�1)
�:�Gd	��P�q�JEaRH�L,��B*E[ؗ����LǏt��\�w Ϛ5k�Y��s�_�̀BbM��慷kN�CX�]�Ō>*����W���3�9��� �ۢ0�o8��g�X�LqMu>���Vdi2$d�g{ڵ�#�019�hM`���5`��J)5�W�0�ug�kz����G�3��j�Yp�~I&������ѿ��Tk�|�ߕ��3���+���Z�c�8p��b�{���#o���4jU��'>,[���@�yn._���5j�~������cG�TM��t�ع*x���&7V���6��jW��E6�P�7�瘗Z-�$tQv�9n<g>�Ju o�)��w��dB.��)�2�߷�-��㞞��+�O)d��ο~`z�wo�����Z�I"�Q�,��l��A]�z�s![�<�$nѝJ�����q$������a�� �`󒘂���aB
b-�Ӷ��$����7�w��� �	�(ܗ8��|�+�>��'��ċ��{D˔����2
$Z>�c��`��q��X�xh�m[`���έ%���Oh����;˜�����9  g�Nک����o��0���]\9սL}
�"\�vI�-#��_	W��s0#��->`���,cNbMHxC59�^��`~�~^s���?S��sgW�ޏ� ��2ѱP�C�q�hs�5�<PK�q�Fu<�g�߇y� �g[����3G�Ŝ�L�ٹyU��X�7��`n5=����!J�K��khQ�v\Wsy�--���٭i�^�6�Ĥ*A�$�_�t�]���[�������\�Հۙs�y*����C����|�K�����%��Z���c��z�j)E^yy�lݺU�����;SR�_ 0v�]VB�yG{F�'8�ɶ!��&G�kU�[]T��<c�%|�3R(�lZ�r��FK�� �\}��g��ʍv�e���+q�J��ߤ+F2����Ӿw��?=6��VG*W�l��I�ҧ sz���$��غ,pQ�G0!1��v��n���EQ�	���W������AT�S���6�h!��wJZ>0E��%
�h�R�s<���s�18$\����-���8+��ҭ߮eX�c>|b����8��6�����-����>���h[0�R�m۟�g�Ɣ�h�s�>)� !�bM�����## ��ar?b�B�����C�.l�v >��d��^���j�%ρ�>-���9��o`����0���984���o @�G��ov��Cig��b�K�]nr�g��s�՞	����gθ�v�q��ǹ|A��`��"�>��Uk-8�릀��B!�̌5�p���#�)�ܪ��_��3��f��k�W��7�6��$��JSV�c.}.>�1���S�����r���r��_��!d+,��P�8tD֮�$3����o�����=;55#����c��ߨ"�j�ў�޾.� �L*�eO�`.UWm�|rIe��1��R�/J�[9|H�\�������/<ObA]���DOO��䂟�& �R�Y1`��K�w~�ֻ�?1���\�F�ALJ.�r�l5m(�é�mjGhc�a	�%Ȕ��X�fǢC2��ݍ��!C   P]ҙ�3p�̲�!�K5i��x���t`	�X����}&cB&�2�u����~�gD1#Q��:K8}����������K�l��i%BJѺ�!�$��z2�Y���fn�ؾ?.�l�kc��-Չ}F���-�� ' �!���.���)����P���d~||L����?�OP�R'ǊW�.���� ����) �eM�l���6��IL��lhx�9`Z��� sęs>���_ ߡ`*�6���),�q�+�0�y#�5�{��#5-Q����|aQ��.���8���3*N���`�>b���ji$� R���[����;Fʞ�OT��C���$�k����z�:��������k�u�9��R\��]6�}r�Ȅ���Kr�����_�'�ƌ��v��L^V����y�ͷ�a?�����K�4B���>4�M�s�I24�/9�D�@{��L��2�(��:� *&��ȓO<'o�}Xf�]h �t6%�zU���J���I<V����iwN���\2uŀ�����{߿�����j=Pu�̑vP3y`����H�J"Gm�2��(5�����y=�?������}<��ͪ�|����Jr>��0��1
t	�V�F�W��z�/2C�l+1[bo��O�b	��V
�3�`���ϴ�6ծFM�gD�Fp�jv�G;����R��3fd�H�}挀��^}�զ�$by��{��!�	b�>C����`�ƞ��{z�C2�sm���j���}��+νf��K�"H��3�I�=H���pz����C'%�����Yw��p-~k�M�0%�}E��m`a�r@���lyԨ���܂�]���?;o�]?��(0'�X*We����ZU�W0Fe*Q:�ęW���\ؾ2a-J��̹��^Ԅ��v$�g��s��|楺Jع�@���_����%��������w���\�����! ���yy�g�S���\|���%�M��R�݅\�ٳ�eٸi��;51�L��c	��1���&Y�n�tt�$��D�R���u���y��s#_�����j�-y�GebbFk}h]�$$�E���+���Q+W�{��+'�G�{z��0�ɽW��;�u�PYU�'�I2�c\�ୣ˰�;.������4f���L�AHU��n��oA��AB����l�gq��!�'29z�MF�X+}[ɏ���{i��!����r��ݿ��7_�9��-	
'!�*jH���d;�$�t�ᵔ�5�)�Q��-2g$� >[��L�8r��cd��:ܟ�������N��>@��; -�����1�$��!����\nt�5�cm͛˿`�+�j�	u@Ұ�ޗՓaC��8j|�3�UĬ�� �]�4p-�-��J�ڗ >0dΜC�,������6M�eh�U��ZuLs��kN���������j�Eϛ��o��=�2d�o�fA�{�X��[o������m[u��V}��=Ǚ'��-��N0W�_��������� G��\:��F ��.�/}Qn����󇞗���,�1>l
fCŚ%�>H�`�;s240(s3���SO���X>tӵ28��D�!�tV������K*�C3��1�����<0Ü��H,�Ɇ�k���$�he`�*�'T�~2�C� �ګ�^i V����bI��r�5W�9g���t�������A0��q��VJ����u�#_����V��@2Yd����;��#�i���.<x��k	�Qp����
ї�|�%�$�V}�yd;Q J�h	.	�U��~��9:>���9��/�F�ɰL��X��{:�Qm���+C��,�����M  H�^\�gdjp/���f�s��W ����h�Ŋ+���V����95���-��� ��(q�x@�EU*�+C��!�_"��(�X�y��e*�K���C�	8��#���7�eM�QӤ��g�� ��p�>���jY�
2*l?�%��3k�WhU���>�a��Y?�D�Y/5��5�P[cϐP;���{����h)S�l�5](�ȑ#r��1m�[��k��F��,na��#>Z��$i�A����R�vuu����	�/Uj�5����kZδT*���y��n�{�{U�~�y��˻��eWt�9^f���ZY�ɘ�:s�f�j)����ǟ�]�+��dh0#�ӣ���+=}]R,�<��>���ؤLLLI����:M�K�Sհ�WKowR��gaZp1�n�\���A{�����C���O��\A��1�|aN��;e�i���W��Ĩ�_��뱎�W��`�ߓ��+���'>����B���:��-��Dq��$$���k1���'�R�<� `$&$x0�F�S���'ƸǪU���wKp��%�A�#3`�� ���*s{>�g��G�Ďmɽqd�?x^o	�΂�={?Ü,���9ֳ��-�O񙌀&:�a���s����c��d�P���G��+����6����L�o�aA�T�=To�ysn� ̬Y1�}*R}�Ir����$�	�1��m�>[�Dd��>�} �@��p��<0BV�c�K�jZ�K��y�s1n��!t�~����̂�_��0�mZf̮��(F׎��������j��M*e���~�G����&=�h�O�^�$T7^g�f�,3�s`��+�$J�	�d�u�����"/�s.M0��u�]]��$�r��o�^�����Ą�wn�]�r	�3J�:K�NH"ېL[ZRmi�T,��{JN߸U��O>+33c�idh�G�m	���_���6�08==+ss�:�y���0�HTUk�q��O5m�*U��q�F��('"ccy��}�پX*������'3IY�j@���B����U�C?�t%��=���[1`~�m����?�R��I ��v���Nbo�ꎯ�KM*Ro����VmL���H��`��+#MP沛�m��'��y�Z��q�>��OT�����d�*U���4%;/��O��/@v<��Qb�^���g�c��α��Q���ӼR��X+UU��c��=�9n���U:��Y�鐈�ö̰A�]�;�x�L����
�av)W��$$��ЛiG�6
��9�M&PY��@�<C����_]�0�Bs�LzM���� lS2�o\32Q����s�e@�w��9[rN)%���=?���}�@m��.��^���v8���9�Qb;T�7��>�5��E��(.z�t�l٦γ�ZYP�!z��8d<��j߁�?n��),����Zuy�5��]5*�Yuy`�3&Ҟ�O�{�|��Tg�G}T�NLhR�2@X����P5��ʒL'$�˸�>my����G��/�T�<�ʪ�A��Y�W_;$�xC2816�`�םdn����@**��θ�rV���U;�\7�QB���6����cR��d~� (�Z���L:.�]t�T*��{��-󅶶`���4���#_s������]�S.�y*�T"�`�Ӹ���s���0S�N�C��+#�+���o�;'���'f�?�vNq0�*��%� .!�FZ#��=���ZC�?�����\p|f�D�O;�(�[�w�)n4�@P���0 �a��{H�L�@ؒ��App���G9��D��  h ~��-����U�5u�q�@�浥��� ]��܃}g�`jB�s��sDO ��Sw.�0Zvu���k
5xHة^=��-�@��;��{����`蛁�֣����Cè�s�Jѥ��8���w�nٹ��Yf`�y����=󥌗���[��ߐS`~l�D��yQ��.�\.�%F�`�Ɖ���Ӣn65T���XX*f#�0�.E.5=���B���V�x���.�h�&�\�H�����%����dD���G>�y���������l=m�LϢ�}]��K�196:.�XU�o�"�cS2;Sh�y��#�ĩ٫���[?,�׶;1.�h���*VM�S�Sש!2=[�C�Fd�X��BQJU�4l�T�jeQv_q�$��������;9O�� ����;��}�����TB�AL%s�y2�h�����H\S���x*A�i�j�'��n��[��`n���r�>��k)���%��(�lڿ�I\��    IDAT��H���%\�� d�"�?>�(`;N~��\����%�8&��0H����ƞή&A�Z��0$� a�E s���.�c^A����6�Zm�='8i�Y�NT���哙3_�qkm5�)� a�5%����tM+F��0�p��a�2s���!��A�jz�?��>�q͹�,j�,���'��,�cA���^u�j�������l7��@ �9g����k�x�U{�s�qq�8�U;ς�!�'��+#��z0�_|���B���
�a>{�������gė�W(٢0	�����k2�a�t��u.B�D�G�\Tt;x�׮�B8��D/ �9c�dsm���!������>,{��#����e��^��OhE���^�UR25>)�zI�>{��L����T�dR��~�Ahi�ʕy�{��muO#$-LӢ{0��k�6��W9p���狂">�T���ZU��낳��=�P���{?מ
^���;�� ���F�7o��?���[+�aFq`5;r��0�vY��in]�T�c�6�.ԛ�CG�\�v���`�܂�:}��H���6��a���T�Y��'+QX0�"�>��lT����I�2:Yf�c�϶�:ۮe����
���X�A+�%�W9$j$H�0 �vL��#b��e��7zM3�'�m�̰F{<��O��u«�@[�ȁ�c��r�k[	
'����\�Z�����~t�����0�)�kׅ}$`sO���9�����،����ޫ�%�^�2��?�Ih��� ��Z����,R��Ѥe>�����?��=v�X�^%����BA3DB��Ƹ}|�eW���"L+����贩r���g���:���6vW#=���g"t� H@��d�S��	B�w��-����$�g��Nȷn� ���47��тX ���A�{�9y��g�ӟ�����#���Ў�-R�h�ŅY9g�)��errZC�ܚY5{ ���m/���7+;�k�r?��m��:��;n������:��· ���%L�r�ygIoo���ξ1�j�s]m����>i������V��o�������"�<�p9�S1�O�f��Dw��+�����(Q2����e�P�&b|b������k�1`��+�+����O ���:�m?)Y���D��ZƎ�2'�Z j �˘'�c ^�ŢJؚ$���r� t��Q��|�vܸ��h�)� y���8�4�p�Q�aZ��$��Ur5�u�ք�����ͩ6UJ�:w�{e������}�� .t�2���k�}p�2�;jZ��Hg��w������KS��O���<ڇ��J�d��yhΩ����z��̕�;���}����Ϸ�z2\+�ٍ�EQ��o4��L& ��u�WIoow_0G��Y��)DY0wH]D�?��������^��fτyI�~G��`BBh#��#�����?��M�*|��]r����ӷI6���b^�I���70$g��CN�����_n���r��ۥX�S�8��#�x�9�`~�9;�R,��P�/��k8��l.&g��^���T��-_%��V��>ǉ���Z��=rB���a��� �o,�Ӷm�5kdz|�Ⱥ��_h�$X	����aEH棣������ͷ��XZb��֎�e1AR�D�6�nl�����V&&��7��y��Iʠ���=���� g��O@Itx�kա���s���:J�Cհ}�}o�yK�ȭ�f��@�`5�!`رZ,�Ŏ�F��-����:���<��� >��� ��Ja�^�äe�@���c��ϸe���Y-O�I�T7��t�ja�Fc��5��p���ίu[8Â%��Rr�HK���΂��>c�<�>�F����*�v�`α�����ݎI�D��?��0B�{�ɄC�"� ����Q�a����,�q�s�s>�|��6��el�Y��7��Lz<��?Ϛk#4��F1LK{�Б0aL����+ޥ���*�L��C3E0g{&YO�ɰ�R9�΍-����[Bk��.<��/]��T����0�OMm���ٱc�twv�5���~��+R��假��rUC�v��
�����w�M7}Hλ�t�T�̐�uIRҲ��C��0%�w�B��OJ��LU���H��Tw��r���b�޹Am�s���~�[{�)���&��9<&33y)W�[S�陙�fzY֯[-�7����鍛�~%��[k��MP��������߾뇇G�w�J�vx#4�%�q9�Cw�-V��%�-"���xSr�l�t��WJ�V"!��O�-��.��jPK�	 l�ZIž� ˽�����>	R+䤥2&Ѳ���Y��q���FtRas�N���f8�Yb�y"�0��C�e$��h������2#Z��|j��d���,��4�a;aF*]�D+�(�����A�k�L��Ɲ$���{׎K����� !�Z�g�
���]:�mM���s�k�Hh��g�ԭ�+U�h��=�y#��I����PM�^:���)�ϣ��+Q);�Q��o2%5��_���3ܣ�����Z����_�9�t�kHF�;������ �"4�Ek8���k������E s�����C8���/C�3�a������<�����>�����_�l٢��������W^�59���g�K/�Pz��%�@�zE~���2S(	*X�<s�F������j���w�����/h�ߙ񊌟�ɉ�����M%UB.�eu~P؋N�n�9��Tk9��-�OޤR�}���B��_��t�H�U���L�S�5���sv����������H�c.a�;�oE���W���[������A�M=$�Ǵj�rЍ�n�'�.ƙ�`�Æ�%�����@K-���;}0'���{*�>
HI@h�#0[@����:PV�a{>C�k�ð2۱϶R۳��i�n_KF��NP�W0���{73�1��U���nE�kՠM�0,{K "q��)ƔI����H����@�y��)��4[�j��- $�p��!�y�#�ϰQ���0�_��$��4n=�c�'�Z�H�� s��|��TX�*Yh8 �dSiY(�р6�=��0g�SI�o�ށ�;��j�,�\N�(G��UA��� [|���DB��� �ҐƑe.��WXu�L��N�ֆ%��^�|W�84�\C���Uo��(�P�����d��|]�0�?���s��޶�؞E�/�;����u6=�;�-�c�\�`�=�{�5j�T�?�} 1"5���+�Lf���7��*��Wf4��`&���9%]�+���}�2(�}���D��M�6�����v9����wI_w�fv˦S����ɹ���uٴa�2���w��3w��k.�x��2пFf�J251�`5{G[V�ZXt��8�U�����<k��r�qu�V�3�9�
[�S������Y��+U�O&�R*��@��s�296����{���!�¯M?WЅ+̟���y�}�[���l�XVH��9$sݼph�E��*��K�˘��}���D�T�z��"1� h���|+�6A{7'2��%:Q��;�>�g�/VZ�����S�W �[J�[���`�Ԏ�6Z�O�	�1=.T��ٍ��f�y����I�8����/���T��F%�K7���:?�*��`���Q�I17��Y��Ŋ&� ��5 NP#�\����#t41�A[p�+4MN�T���xa8l��LZmυ��&5�АNH�`ࠄ��5��,�3���yIg3��v�ߡZ���	0`\�7��ӨIp��%
H  �A�f$s�OJ���TFAU��sjUP���b`�:�:����.?��x���1�n��?�Q��	{�r n�el�Ʉ$<�2f�V
�	���h������˯T��7��mݥzen|�=��p�
��!�� ;D��B����s��;@�M]�*�������_�,u���nX/�=��ڗ���y�g�i�p|���]�f�_b��tw�c�?)o���Z#.��{圝g˭��*���5�]*}�(�H6�&'*
��#r�雥��C��f���=�C��FI*�y9�����j�c
h�R3�6��Y
qa��ȱ�Y91>��P�c�`�����Cv]x�L�OHo_�7�������ѿvWV��≽����?������F���)�D�4�E�y3��L
�q4�QmA9vϛ�$�6�\H`<����@�܌FI���@|��g�>a!���`I�ҹ�I�x?����>�}��^k9^��m2􅟣��@>��a����� *��e�jkփ���@�7<=ީf�#ד́�K�2���� �RrR�0��ٰ0 �j  ����C��2 +e~jN-P���U��!h\p��ش��-0�F �lZ�9�aL!xb\��%���7�R}:�4)�a}�x�p1o8�ׂ�A��G�T��Z�f@��K� c�t&T����Ήz%�~���%u|S�vP<� ��\9��|��~E���3�������g�2��po5�E��b��ͽ��r+��C�Dm�>�T�Lv�HmՍ0�u��̱7�7d-s�/s�u����w`�n�3�˙��g���?���)-����{s��������������lX�V.��ٶi�fe���ǟxJ�S����N���]��o|K:;��z���Hww�D��.��ԬLN�M��h2��w̌�؏�*&|��W���Z��Ӷ����l�u�����X:�9����c'
r��X̱7�V*��ё�K/�%3�S�љ�I�����A� �w�ߊ �|�Ɵ����g�յFBҙ�d��j�I�������K�O0��[	4�����u���FBOX_��!� ��n	���q�����21��Ϧ�R*�JT{�������gf,3B����h�d�	n�.�o>�555���w�'Y{�L/w�$>��J�FA/�)W�/���-�r��� ��1	Zy � .����T� )�7�͆���9	��~5�)�<�U
M&U}L3�~��R�$ߤ+
Q,���(z�s �/(�Ѷj@K� VC��1��c�g�זJ�9̍�0?o�X�V�>Q��8��A?� e��fW|�Y�B�9�> x£'�)��*��?@ݽ�Nb=]݂:�]�ʨ�%T�C�lj{~��i��g�侔nA��{۞�-F>�w��Z��t� X���g�u��y�:l�kbj���Xת��;30��9�U�X_ͥ���8���������Z=��9�/�n���i9|dT���n�M���Ȇu���Ζ۶H�Q���>���K������:��+/�[�{�tue��I�����DUF��i�����f�l޼A&ǧdn�)�t]�	$���P��e��!Y��SD��|0w%��r��5P� 2�S�2r���ّ�vs�Z�.�U�/S��t6�`o{ח����;�WJ���y����(���A�9�1�K*�������T͎_���H��dn�)<5K<i�R�[	��d{_[���S=h%��Y��:¨}1�����e8��:�͐�0�����U���{�c���2AH�a�sI;*��Ç�����e�T�~�FFF���*�C���~���󟕴8��+��D�G*8CU�q�Ǐ+�ezL�F��Ƶ�2V�U=��ѦT��2�s��2���RT�\Tr�V���@��c?�T�x�����sf3�X%�iu6Y�t�5����u��q����l�������	������{����Zq5��a�5fE�mY�#5CK����M�5� ��\���m�D0���?$/i��ڏ�ëd�j��q>���e2BU5��E� cR�̰��	�d ��� ,Ք�� ovW���c<�����ϗZ��pLUI��jwt}�Z��V�_\��#@�0�"���~�wX7��9\g�����G?$��?W��ۧ�j�tF���}�M��W�V��^ٻ�5ٺy�lݶQ�o�(�[�fX>*O>�*ɵ���+����S����?����p�k�����_�Ņ����d`�K�o�$'NLI~�sTeb������n]O̩fw�3��z��Ձ9$��|Y9�·����NԥR^�{�U2?;'�D㉡��ϿS�����{?~��>��?,��\���L�M�m�ձ'���՜���1��J�V
s���ͫte�U�Z��^C���[��Q��r`��|5;�E�R�r�%T~?�NT�����gQ��*��E=(T�\N��(-8��СCZ���7��ձ*$Vt�Ґ�0�̞={�`���֕ g���`9�TY��E��>� ���f2��6���$�9�p�6^*V�;�z���w�+biT�h#�ɩ��R��t�Rp��s ט��}6U����t�T���VkL~&�V�9x=SI��h�� ���rϡ���Bbς*X;�3�;*�`�g@=�5��h��tF����XXP �8��}����*p�V �����RJ<Z�X`��>�O�_[G��%����o��ڞ�Ɇ��dݚ�����	�h�v�r.�]B,��,s��t�3��>�o#)p��g��1�������7o�K.�D���=�`rzJ�\r9�#��!2#reP��Mf�PȫV��`��-�"C����߳[���je ������ɧ����뿖'J�~�q9m�VY�nX�ܱU�����&������bɃ�r����Ǟ�����|�T��G����tM
�E�������s�69>:�`ޢ��O�reNV��M�N���5�H�(�ȝ���B]:����.�-���\��0%7�x�,�K�������S���>���y�ш�{����~�?U�A�ވI6���<&Fͮ|v�вb��.T��W�\�LVAI�&���/Ջ�-��z������b�~Vjf�-@�\5���o�=�D���J�VB�ڪ-�?�l��C5o | 
�\(����^��U.��XA�F��J׶o���>P��N;M�Ǝ���y?�$��s�kԕ�;.�P8 	}R�0l�锤2I��"��_�q�LMO�k{_W�tbj\���ծTe�H�:�L'�.5�5l��3?�lù��u����V��YW�z&����~Ch/ ��O D���/.�Z��ɩ)y饗�Y��w\w�ʞ^Pg$d����c�ЗM����;v�#4`F֭[�����駟���q�©����9b����W^!c�� �:�;\N��Η�z@&�ƥ#ۦ�5���b�o| 9�z���������6�P������a �r�3�I�5S���3Gf�L_s�{�������T�-w�%���o�?�{�`�q�f���˕vACA-�E�)T1� yh�������sDE�U�9��Û�sFx@�~����ݠ���5;ڡ�#��C����/�J^xa���}�}�Y�jP�?w���"}�]20�Y� ����뮑�}F�'_��HggZk�;:-s���e�<!�mr��[�����S���9ՕB�G���P�l�J0���K�>pK�<�
�n'R)��QX�\74L���Ԩ��}���|^����>��<�N o��+�3��/w���ϼ�W5��'%��J�=�\T��jY�m��8�d=�&���I��(��R	b�4n��H� Gp��'�jp��j�fm��p�`0^h&�(��Û�&�ސ1���JԶ�V#��P}�{���9�L		��@U]�cm�0C	m�F��ּ�yT�s�K�&�P �mؤӍҜ�7�xC `�9�X�sL�lK�s�$���j� m?��S29=�j���B̐g�S�LZ*����H�<�li���~�̗
�ޖS�xg��:�9zxD^�U�%S�?0 s��VD�L]���]��f��=,������L���oX�o�"O>����%s9���K�� �Wi�v��{��k߭q� Ϊ�T�=�^'o��W��%$��h~�䪆�*(�ē)�y��
��>���k��햛>�!9q|T^~�y�W��- k��XC*pB�R(�ӷ˖��    IDATm�塇���k���]�l�(O>�������|A2mY�/.J<�Q���Ԍ\v��2~bL�>���wH��׮S0WM	����	�rp�	ܖy�Yṥ
�F��2�~����酼6)m������
���Ͻ��r��kuLE�+���ΰ44�>�����S�
�9"QK�^���w������I2�TF3� `������e�ֵ�{�w��tڑz]>$�=�G��Ͼ"�>��{�}��-�fxH�n\/���І���{�j=P��+���o��_yV��/�P�Pw�.��r�XI�1����L.)g�\'s��LM�H���%Sf(�<��a5�e9��Uj���J����ƮfV��
��'"�$"�"�����\A���i�8܍yK�{�n��ꐙ����]_���>����7����F�-?���~~ϿS�X\U���v] uBB��s�B�g%�UY���`c����K��u���Т Ŷ�6����͸�&�m\� ���C1��$XZF�����c��m��K�|F��Ѭ��=��4 �{�6�o[�#�7�$Xe#6Uf��	���g�pB��I�9�=����-G�AF*ՒƊ��g��W_�|�Ղζ����|M�J�T����X*-]=ݺF�ΜL/�ʍ~�<��/e��1iH�����&)���w�+�XR�{{��T��]q��aiK��u�o�w}�F����u�&�H��ղah�<t��r�gH=���i�<6��e*�7�j�X\�y����3O)(��V.���]+/<�lX�V�@F�r��"�,b��d�歲f�:y�_J<��1|��=tPF��tV������ez~FH�Җ��jY���]���]~|�]�2��l�ʮsϑ�^|Qj��=pH:��Z8�9H�A2%���cq9����}P��*ʶ-[\1�X\�	��9���w߄bώ�-�lϮeԹ�� �5���J%�Plm ��:`>wvw��W_-�33@��nȼ�j��dN0������XB
s-�. s0=�Z���O5!���yq1/����>�)eO�=��G�������/��w߫Z���ٰf�����l(�������yP��%�ٙ	y���k_��20�.�zQ�s%9q�(ss"���񆜻k��� ��kˆt����\�w�f�y�I[6.�OT� �\i��{�N�!�j�����t����I���o��B�$�xC�x��}��g.SS��W������������o.���5�o�֏���_�(���۲���T��!��+͂>��A4�,�s�
�@j������_gu,�X�c?�{n�ZS����0��%Fl��`�$6V�o�h	�ܟ�v�d��9)j8�F/�S�9.�Um�(��� � �V�[��'���5�a;���u��l����1M��z!W5���oɡ��R�:�o"�Ν;啗_v�e���b�7�D �f{o�����r�G? /����NO�uӳ�����}v�xe��|V	2�rKdU������̤toX-��埾�uM^��r֚��s�6y�w�Ż.����Q��PPB�o��V�X(W�o�y�٬۲R����o�Q^x�iٸv�~�m�jf��K �^�Q�ggeh�ٸu��}�ݒ�lW��{��7}����@�-�7Jg{�K:rlT�1�#'Ƥ��Wv]v�|������]NۼI޳{�<��CR�����<b�4�R^�='�TJf���!ٸm����+ҙssP͟{�92�ۧ{/��6��ʔ�M��������'V�c���q�]�)�<�<v|L����;=�&W]u�$�	�w��!��QE0���4�0�`�g.�/*��\��u;&�~�V($�� � l����+2v���i���rI��yEn��}���oȭ�~_�=�|ټq�z�wd3������~@ˋ":Y������G_���q���R��d�hA�'��0_��bAv]�UK2=�����ᖞ�y��>g�^�Lo��QC�@�$@ z�b�1n�َq�8qcC.;q�8��Mq�$#��B�PA����sv/�����>k��ᳯ��+��f�.oy��YϺW_˨�m0o��m0��l0��|.�={ף��9���`�NI;V)��`n�^����-Y5�r�f��}�q�?�l�9��O[X�n�����������cN:��^��7_���?�ī�T�Jf��P1���]�6��D��H;��^ڔ�8h�A������%%{��k���3a����E b,ߩ��+�ו����|�I�q�	�5s/�xbչ�4��mL���x<�%�Kc� fc9n�ʔ���(7���g�y�L�������&�~�g�����6�x���M������g��{�����z@�lj����G.�c�x�/��=��>��4���K��g��}.z�C48}��@�ˢ(��|��p۽w�w^�����e���Աkx�޶���Ul3?2��L;L��a���>6�+��|�ƛ�j���lx�[߂���f���`N���z6��M�19?��[�a�Ν��m�Z��L/?�\�윳Г�alh׍�6��|+��J�T��o~߽��{�+��݈��"2�$vn݂_��*	l]7�˾2*��B����q� 217������7���w�mG�TC6������� ��z{��70��C��#0��^�=�  �U1of�4NnE0����5+����I��/Fw�;J��*j��B.tp�/����ô��~�"�[��
�Y0<�T6�G�5,���xj���`ӆ~��/�/<�,�mۂ��^;���k�y�9�s�>�����;�<k��ە��+YV'�eq��������s;�{
��ֿ��..�삨_}%=��r����Y��/A�^��T�	V�҄�<�nb��M`�|�x���2���=�:�>t5�ߙ�eLM΢\b�*kE0�����^��=;p��/��#�ʣ�C�qt��#?k@��I�瞛�z�o��g�9�Em0�*��R(
��G�(v�D x�]�?w��N ������NLB�[<c8�4(�i3�3����fp�OZ������ъƻ�)\S�h<�����~�:�i\�/-�0�5��<�A�Xcf��]�k|zΏ
�м�t5;���8G��k��$X�9Ό����h��x~���|��1?=e̊`�K�, �\�R�4�+%\w���-��O���h1g���+w��מ�r�����`c��_G��Dw��\-��������p�{߅k��3�v!���x˅?���,F{Л� 'jY���	���o�+7݌�^un��f,.�Fy�M���7`�� Fz��Mj+�A2�|]�>ku����ʍ�`ra��n���f�U-a�������-l��tQ�)G5�Y��u�{r��]௯������u�!��B>���u��׿�~��bX-"��qȐ	t��f{
��ſ@~p�F߽�n�r4+5dI�?���4m�knY�Q�s�]O?�{��c:$���.�M�uY��z�s�~��Y�̋Q�5�/���`�! -�X5\Q�{�3�=�X��,0]$��_o��~�OS`b�c�T�Y 6��5�(������	�{��2+('����,z�pɫ/�_}�q��/��Sw1ت��Z-�����gqtb�ܽ�w��3����?��\r^�+�hV͟?9Y�ѣK�f`���Y ���<VW�P�c����=�̓�Nݵ	�����&��-��� =�A�h��ϗ0~l*�t��4����:���~\r�8r�hkp��S���֋�>�I���:�����K�8x�V$��B9G���R}45F)*k)0��ٸ�v��=�9=h�,�A�K�^� <Nbq-_���3��	���2��pM)��?������u�O�*���iN<#�:4�2蚪���� d�����X_␊�k�5�{��O?�t3������Į{�Z�L��M�J]�j����G���]#� ��z�_�����D��@�R2f���VW:��Ss����.����q����s�:UF�	\��\|ڙx��]H���;�Nbia�6m�r��'������x�Uo�����==H6�)���K^��lކ$��Q��V�c>��a���s��������]t����MS�� ��^��~���.�&Н��^��k�$�4�>�ſ�S`�K_�o�{�)t�U�b��1���Wb��1ԗWLa��ֺRk�h?�����i\��7�˷ފj�a��u�(.<�l����"���Z��*
�!�����$����������$��{�i��y�t'�������`o����7�-כ�� Tя���B|���u=}\���U����}��WJ��5m��p�*�j(���P��{D����\�lrb�Z�x�	?������`ш2La����b�D��*~�w~�ӓغu3�m�b׹��/Y�w_u>���q�Yg[����,f�'1q�0;��ժՑ�u����7]�O~����/�e��G"�X�_��b�338�]���c��,V��hF��8��[�̛�N9u#FGC��&���BEǊR��5S�k���*��0g�&��������u����a���_z1�g?�`��G���n����Ng�#i{{��Ax0�<F�&7�(�Q��ރ1�UИ׌=8	�|���O�8��Ϻ�g&��m�2�fo3�'�4u\q�#�q���gN����l�r����mY�� qa�k?���� � a�9�y�;3��yT�S�k�h�~cccv,ӡ,�<6�m��z���RVMV�b��z�f?y�qL�΄��V�����ށK_u1zs���#��`���r�z� ����v��|�䀇�yiw#��w��K�6�;v!Ӫ�ڬ�XYՌQ���=�(>y��qٻކG�}
�=�)T�Vp�g�m�Q^X@ww��W��9�G*߅L��=?�C�=���p�XHa���(�s8g�i���Н
�~me	��0�~�ZG�Af�n|�����c���}rv�D�d�GFp����;�3kD�|�ӁZ+������C���klػ�8�f��z�I��}'�yӛ1�ɡ^ZF+�0�+ڑ9/.Qn����_��m(��_-�I\��7�sOۇ�T���͢B�2�Y��z2�r���=���H�����(.DB����������^.����WW,5mt`$4���K0_\��%D(��4-S��A��0����d*4JYZ��Ј��t�����-�m��V��~��9f�'Q�qƾ�-���[n��������/\w��Plhnf��VCZ2�C�������xՅ��W�|=^��3�^Oϓ�X�mf��C��1=;�S�l������by)�yا	+�DK��Zu;Oـ��m��ە��W�������m��r���ւ`�V>�7�X^Y��W��s���os�Ͽ볟t0���^��n�~|rzM��4�*����ԞX֕��m.FNZ�� �l�#f��XO%4�4�%rk����d2�߰����q���4�X�̂kŢ@0��o{��׆�sJ��9.i!k�Ú+�kJ����}P�g��i�5Uz~1T��@X�Ƀ7����7�RӼu@LV+�g$��{��-e����j�l)���\�*�5Q�W�i�%�?�ԓ82~���l:�t��_��w�]o}���h�U#�Ӆ��>���_\w-��1�ka���,=9���v��󷜂3�lE�\A�7ԟ�i����	��Ñ�)����K/�G���b�Q$���KNن��E3�QmXjS�-z��bzy	&&�T.[ ��=x�%a�p/jKed)>T�f�Hu����a���xO>�F2����P1��@w�8��ؾn�>�ҸnQ��L�4��805����O`�����(�B��L��37o���;��j6�Z_F�R�`���`����⫷ݎ�}�3X�j��a�Xj	��a��y��BO�+���ꛋN=�k�H���= ���Q�q0�o��R(5�0[�
�Mc�k!�6�%���1Q�<��if_ZZn��q�
��k��m�˕b�d�����FF��c���f�B:ES{��*��7[����,v����o~�;��[�Yg��cO<�R�]�*v�z0���H��۲F@�+���^���{�m�(~����Y
M�3Ncq���Gm�nݱ�6���yKk4BED+��̫�e�ع6�zv`�(��ʹZ�d"�9��Q�`�}��?�Y�����7�XZ"��56:��B!A�z�t0�Ʒ�ڛo��g&&�7���H�\�%+C����� �7�5sӜ�aC	0�1�|hEy��N��"<GR�6;	TeJ�6fج>7��z�^��o��@*�W�i���(D�*5z�f`f�`��{`���5Wv|��5k��[��7�]���4j�x�����i>z�W#��1�&5��:���}�A��`F���r����	6�ʹ�l�(`7��|���g�4�3d��F������!�h�;� �*�t������<
���2Ȧ�'�
821��B?��E��>���<�z�H2��i��}8�6\v�y@��j+���T����E�\Coo?�NN���|�7������snz��mC�Tľ��P+�j^�$�ni2l��Jp��O�K7�Vo�&Zk @�K��_y�{�g�VԖW1�[��Vծx�s���߽���WQ40���Wq��߁��?��3X7ԏ��l�Qkb�XF3��|��?���1ϖ�]4���B2��D���`cWҭ��rf�m�ط�ۚcdzz̿v�X���'�V��g��Xa �j}�T@��k�z��v�=G��y��
����XV�R=蛟ڄٵZ��	�Q�R�-.�XQ%j�fN�V,Ps���A����|�4����!��>v�x?�;e�0�c�\� Jr'��9K�2������A-���t�,8;=����N��ƀ��[6���..xŅ(Wx����<��Y�)�7ۣ�p�ˇ ���n��Н���Aw7��*���f�$S�,���i�m����N�B����"A��U"�f�J��bp(�={֛ϼ-4��8���Ɲ���JO�F�R7k6�� ��8��/}��"��҃[6��+�O<��B���_���}Ƿ������ %�\�co�̠����ź��6ʴ�`>�BP��s�즴Ap<���a�;[�_Ҷ6N\�����Ƀ�@S��D�)ą����%gi���KE��k��]�͠�������I"��wC���&�Dfv��/�9�5}�n	D������A�W�!3��4��jl �{̮S	G��% ����5?]e涒�����}�Gѕg��.}�E���^��\
cC�Pȶ�M�K��Y���0�M��}쿡>6��,$�Ȧ��60�Tǫv���]q%��N>��ߴH5*b���?>�Y�ܻ�lF�`�R]����ܳ��5W��ƗA´�n��
z�&��,~��3���D���<}�-+����X��ͯ�;7o� ����­
"�����Ҹ��ȓOa�~�Lh�:�Ӌ�|;׏�ݻ�C�l��hZ�Q3!�1������vL�X���f�\�R�����c]](.γ��E!_0�j�TC��7��M|��� 6� #�7�C��Dw���-����= ����wO�<G`��':�>��k�G��ý�� ��d�Y ��Vˁ�i�&�o۸5(��fN�*p,;Z	)i'�f��-[7"Ϭ�z�zp�Ѭ�J����Ϙ﻿ o}�[��f���4-������c�);�k�N,/͡�����I����Ng���]x��Q�,�Bg�Z�d7���1����'����[��b�� ��3%LLL��ha׮��e�E4������h�3��{���jX<с�q�Ͳ`,�Հ��>zd�R٢�u�(YL�����ӏ����Ć��W��$��`����n�����=���\`UV#�1
�mBo��� �]�oM[SD�4Y�I��������]gxeT���2��Ci��w#`�ft�s9�hnT[�v    IDAT/xm<� ⟽�ۃ�m�H���FR�dz���Ō�L�ͤ�(\ϴ���	K��p��m�Ax�|�W��9w�z�=ǨFVi��5-���.��V~�1N��0
z!Ѝ��8���:\3�#Yr���Y/gg	���?�ɳ��(�^C*r~��2r�^q�~|�WއT�j3��&���B�u��]/.�/��7X��H��ZO��ڃ�z�Wp����o�չe��]�ɣ\�ZX���h��|���_y!�mڀ#�㦯݈]���3Nۋ�.��Ҳi9}�Ka_�yڽx��a<w�0z���Z-cn~�|�,,�j4p���ul奥v\J�s��陬���z� �;|���7����^��Ã�ʰs�Ft1تUG*����&���o�����y|�s��s��64@i?�ְ{�F���Wc���i��LNC_��iM��>��;�oFߺ1K��f��/����#�H�'J�&��#����6���_�����A�z�_\� ��.ը��c�
o|�`�9�c�imlQ _[3g��r���+�eA0ޔ���Ϯ~'֍Y59
�&�&2XY-ế���>d����G�}�n��������a��s�9/<�4j�"���/�寂�z7�r�z� �KV�=ס����(5n���#C����у/���g�ۿ�kطo��q���|�j�Ss�5j8��혞��2�z=rS$X�G��5�����hmMۅ¤�q'�r27,���.l��8�����f#4@
(K�}�Ns]-,�ذn���e~�����~�I5��.��_��_~�����j�LY`.�<H��0�˞���Xt�\6&of�\�]�R}�y]����<փ��¼1��<���C���̃�t����M}҂;������~
T���e1h)ʇ�򌫭��b\$p��n�Kϡ�z 7@ȿA �L2��2@�cn,����L�%��y=�3�M 4!���������ԲM���̭ow�nfD5�ge2��z�d�4�K�R	S�N� ��:V�#��4=kwZ+���++˘�<�F��3������O'�l֑̈́�*�b��U,;����}��(p���z!���51Rl�;�����&�V[h�Y:�n�cXhE�X'g����3����0>�ɿ��s��;�����`�0F�[�4�]�Z���E��Q����js�6�=]yT�
I$1��c���
kћ4k�=�Y<w����al�F�{V8fǶ����p��_�_����z{2�2U��ѝ%q�!��?��_b���F�L������9{����y5v������4ڈ��Zs
���w�oo�	;�����	���^$�-dٿ!�Cie��Ǯ�,��D���u镴"��\=^h����1]?�U�E{�� �?=3�s~.�K8�쳱{�)��+�ǖ�&�/}��F�g��)07>�N`�)���(�ݨ�����"p×n��n��Z���H*��d%�H�G��O<�W�|?�fǑL40q�����������㩧_��B���[`�Y����º�a�z��� ߇���_��=��ӗ	��Vk����s�lϝ��X�c��,jfN�K�	/�����j	]`����-�4��� `D���rA���q�%]W-=���-��ic߶m��g֭�š��-'���8�`���������п)��6���ni/�ȭ���E	�+A��%�Z}���Lo�H`��<� C@P�u�R0�7�y�<n���{��K�^s6bt=���j�2#�k��|Xq�:.xx�&�d+������1�����G���8���H��F`f�M�|mذ�4m�9׎�V�5q�#��|�r��	?����3{�>2����:�4ْ���emP�?�b��Mx�{�cf�f�b<>{:�E���t.��f����_1�wʽ9�/��\�	�\����p��sQ�1��"{+����x�r�}�}���������/���vm�d�߬� r�{7M�4*���'�ͱ�p7�;��YPE's��}��[@�u߻�X*2��B��O<s������s�R*��;�ĕW�����I�y�K0Г��Z,J���"�$Y�)�g��>�)�9�L��g����}����;w`�P0��>�j����|P�\-����O�g���X�o�O��@.�F6�2��<�*|Zg/��2w"�4"�x�n�2��^`������\����1��fv~�Ϝ��/ٽ��)���qM�f�����n����ڀ?��ߴ�1�%�TTXki��/�f�����#��ǰek�2�yт�}~������W_�L�1+8t� ���w �I����>�i�/� �q�x0y��B[��JZu���~�*�����~���o�Nc�n�Gr��߻w'��:&&�P5�����3'�o��Hg���B�f;l#�M[C>�;�{�v�-��ĂE�ӫĿ���q� kF�v�.�t]�ݡ�����Xz�?�`>=����-���{�}��b�65�����k�B��ݨ\�d sV�R����+ �������^�-���D QcK�H&m�i���~=�jc���(���2c1�ݛ��̅�F�	<��\<���1^#�=�Qǅ18�0�9[�0�WY���}��C��M3�|�s���|Q�k������[��t��	�Z3�'�1Y^B7�`ʉk�m(*��f*|e��(��%�T�h�k��9g����>�_�d0a&i�&��񥿿�[7b5+�j��p��z$�J��F�53��iZZ�|��@���l�B.��~��c�.v���r�GQ/��_lT�f�I!�<c%
?���	���4֪��h*��8��l��w�\Ş��8:1��� ��捛�T�@+F�׊ekeJ.Ɇ/6�iVp+��l����T�T�Z_�L&ߝI#���۱�
�.f����W���#���-�z��P@K�֚����-��<W=��I{�t&AP´�U$ �$��Ե����S�t�`%
B���	��f�z̷m�f`N�C0WkY��9��=,��c�{��ө&6������Gww�Pw�^�f+������܉��e�����3�P(�������C+x���g�6�,謌g�z
?w٥ؾ}��z?~��'1;�$�(*0�[����ϴ�a��LP�������z.��lz�M�*�'{��S/]�ڵ�^+_[.����5�� G0� �d	�woF��&ȵ��p���&�Vm
�bjj��pM�3�^X^Y���Ǿ}{1?7S�������$���������
拋���~񖿼^U�� Bȡ>n�RQ�� 恀C�#����K�Kf��t�υb�G���a�1	��~��=���n����}l^G~i�>,ڄEf�w	bj3� J,GU�S��g4�4^��x�����f��?�_/�����"��G��	32{��Y&z��2���D��y"�c��J���s�a�3��Z�ޫ���S��fĠY/cfO[G�:pV F��	��9��m�E�/�O��L��g��T�Ճ���.O|��_�
��R���pS����Vzp���zZ3@�Z,a���V��̄@$6La&�a=�-��!��N˾��*������̣R���<Vˡ�<��s_�;�Z)����I�Z�����2����D:��v�B�`�(���,��1�vMU2e�����g3�<�1˅y�V���ػ��bb{�	l�<�Khl����-�,�3i�٨5��_�
���fv/L8LӞ_������X������S����4�V ��Jpˡ�;}�eY�R�`ǖA���(���/m�G�	L�.㮻��w���}�9|�#�3��f�u�R��b	S3->:���<r���-}�g����pι��o<��zǎN[�a��_�̙���$�M50�n����Jg�����+�x~��� �b���h.�صX	�Sv���G�N�X��4�V��y�m��i惃�m0�>+Q$û|��UT�`>>>o{ �bS��+�WQ�UŎ�{w[��������D"���뤂��Jk�����<���^�j�50�fk�D�R(B��9ps�������͠��L�,[ a����1j��H/�DL-��������1-@�	l���f�q�����G>m]C�-3���t#[���	�d�Zc:�����]G��s�#�@�n.[T��[CL�b�f�'- �ǓA�����u��4�Rqm?���t��Hl���*w)��ߋ�kS4��B0OԵ�_�t^��ɔY��c�U���4Ka2o>v�e�#��/�4�m��!��F�d�� �,�B>��t,L�P,3'9cZ;i�q	,�T.��e��B7�K �6���[ '}�� 0�?�ɔ$��B�w�"��ao��R+�J�Q隭�r�Y�r�9��%��:S�2�0fj�i�듡�iw�Г�?N����SjAlk�kѽa��
���K[P k��qӚ�P � ��a���������+��\���o��5�������#n�����Qm������yZ��;�숟�� ! 7ek��J�.<�p/�5�Q���,>��?ö-���ڠ�NϬ≧�ŝwރ�x�Gƙgn�і�MKu�-&���q,�Oİ�<�g�~�y�kp�y;p����<h�4��I�~�����͑�!����C�ߏW��ex�k���@��maaK��u+ݻo�N3y92��*��T��i�K&�G���Ɗi���s���筽q3�*� ���3y*�E.���)��X�ک�����,zzs7����?�Hs݋�uR���lq�g?{�O>}�b�����\�tА��Ө�!�xL�Ĕj&s2��l���=�|�\<2nH^��7�T��7fJ_9�Í&0� �u��uS��f&t1i����M�)��,�3�-{�V����(����˧h�5
"��4�1����i�Z��z�� �b���eQ���P��[D<3����\I��3H����7bˮ��f�3���źT��|vyS���WN����&v3�֐kon3?��`4����]�Z�e:gf{������c����iD�(�[�Z�Ӏ7+K�c�6�C��3`�ǐa�%�r.x�+����Y%B|���xXW/
$3�LV�)7$E~��y�P�94�ɴ�u��C�O����h�.�@U�p� �j�5^�PW�a9jM��mC��y�f\p�v]Zex=	����C���x �܁x,j��f	ݹ*>��O`�M��m����NZ�;<���q���G���b��a�z�J�ƧVq��$ʫe�U���bvz׼�j��������Ý߿�Sv<��!���,�KJNg�����:�??t�}8��=����cl�Ϟwq~	�\�f-a��1z28|x+K5�ҡ!�.HS&��o���Z	[����M=Q^-��I�t uE[���
��e�X�_�H�l�(3|iY+���l��@�t�n�06xM"�X~��x��'s�'v~�s����sGΣ�Ib�e�-�b�Df������+� <����c�lZ�)��hF�op�NI0Je"��y<���g�q�!�(f�����[��-�)-�3�N���y@��[ה�[�b$�*U��s�iz&�A�# �3��5i��a�/(�мj��]��K��g��/0�u� ��ј_/`�AP���k����s$����"z/����FV� ����NB��Q�������8� M㏄ы���Ӡ�#bB�/���5&��(Dƃ�����w	�zV����'h���ב��2��Gt�q��6D��.�Fs^��r����\������_���@����5�*���ɝV�АG̛�2Z�%�ٟ�	.���s�es����7q��Xv;
~���i{�bq����Y��OM-�ȱ)�Vʖ���r)\����+_��~���}��\�J�f�hVbm�O6��t����Q��<�Ѓ�w�N��c�h�ŖLML#�b�$�q-�Ynz7����R)�y3�d:XE(ఇ}2�l��e�(�l+��P��q�u���g�#c2��U92�L��R&,���(���b�h�����_�H$N&>�c�}R���f�~ắ�����3��#��N��v�[�Ɏs1.��c<T�3O1K��<&FC]�3�1H?񺾘��=3��|un�y�Zq��>�t����8(�*��� O���_�ȵH�H3�1��6v��Z�t���3e�S|<�\"���C��Ӏ���Z�U�D�������qaL��k�5��B�t>i��5�Ϣ�O��;�=.t��X���{�ԃ�_�F�z�=96+hU�ӽ�Fq�Ǳ0M'�mk��5ˏ'��9&�����]:����®�V�} 0g8��4>�-�{�~�2��Ԍ�3�|dd_x�ݺ�.`Q���M/�.k�Z(��
.F3��l-D���ض	��v��]��l��d
��^=tԲ�^|��ކ�6����}*�:��V,�T�����Kسw�;�,��M��C?:�{������J�:�<��2	�3��i�10��Ɩ-����o�H��B��	d���jU�������#3�5S`I�_:��Y\D�7��������[��n
�^���:07�"�*�`a�!����!�Tz{X]�b��|ǆ��{���,����O*�����3����/<2}'��uOO���(f�A���� ��i�
�Y2�����k�12{J[���38�׌�`$`�Ҽ�B���k���@����ۉ�).���=�ۼG��Pgb^�����M�,�}_gf���9�݃x�̮y��80o��牙z+G�
��t�������֟���&�G�O���ȧ����Q�P={\(���9��㚴h�_K��ӄD����:>&�&��H`�ï�
�r��`�9e��8����h7�ڣ�w]���W����{A=��Y��M��8}�s�1�����B<F-�ӭ�1-.,��v�ee�Ӻ�iL��]�����Z`]w��tT�'�Ь�=tp�P+�:nؼ	]ٜel4�M��-P�vy0ȑAj\x��8��M���C���19����"�5ƗPѢ|΢Qi3����L���#?BO��;��%�nx�t�Y�����2zz��m��[���E�ӟM0�t4:��kPA�`d���^��e7��ltr\��'�U�Yl�RB��0K�P�j�b�R�������cÆ�����L����,~R���>��/��u��͜jRx.�B���fv�#�u���i��nўQQ�8K�����/mJ���Ơ"��dvs�8�f��k;bl^��kxq0�@sϘu��Z�	�"&(b�������;��͌b`bjq��KL-�,���v�������?�B'-_s��~�$�I���&f�?�����kx �*������8s�q�0:���t_Η�U&l�����Ik��B��G?N��D�q�$N��/<s��<
8�h��5S���(�ym��<�y�1H8�sj��{F��W��ǋh����x�A��}�CL���9��ɤ�53͏R���q��x�m�RCTǞZ���$���`b'X����եvP)30������F��$����[��P	��(j��D3�#�H[��z��/z^��p����3Gp�����J��Cq�|�^�ͦ�H6L8aY�|O=�8Z�~�W���pF{p����
ݽ��+�r�)�09����e�#�[&S�i���u�U��r�{�&ˉ�h�X�V�g�xk��`V��G��X���jfv��gf,�2�fa�:������S��_OO���"h�hL'̿��3��ʗo�����V�\w�{S´�Jx����Ѣ��̴*wh�>�(����y]ik�0�mtt��r�e��@.F$&虡Q���iRq��fP�A�AzM��ּ��1z�,F.3�Rs�8Jq&�6�G�,1uZZ��F�1t��s�:Gs���㙹˸f��5-/dt;O�ƉhE~e��h� h�D/�����~M5w�g�������N�h\МK��H�׳�����2M�_��/�B0�ӵ>��@���{A&~�����A,p    IDAT���p���hv�g�X|Ǌc,�J���v�����r��f�W�0hY���GM3g}����&�׊�P��)]��,���s��,���w����QO�V�
%�*�8����w����	/
Ee��H ��<2�Ӓ�y�U���Q��p��,/L���P_G�̛0��:s�J޽kfg��g�y:ŔD��A�SKS�V]�$�����S3�]U:���� �<*�� �l:��b݂����1>>���P@&XE"Y�Yg����g���3O��C�Ģ�ȋ��I�;��țn��;���^Z�N@]]y�7E����*�ԣV��r���Q�$v�$onF1F+����(�iifn�:%�Q�c'@��o`
��Ǚ��%0�@�����V������៯�9��d�,� �,E�ѹT,�ӕ��k�޼��
̍�E�|�L�_���N�=h��u
�����^�$ ���}'���t�\:Nc��N=��VĵPO7q���ょ��8Ӓ*Z��j,���<}���{o�2KN����%�B�V�zi�4�^P�w^��3i��W��{��{W���ә���o*���z����拼벟�Ԕ��k�̇>x�y�\A��v}�+���x%����yYB�O#��]�}$�ˎo���D+�N1[�a��J���L���m��������1�]Ys��Qk� ���������QL��/��;�~l������:�9[(WKf�?��1,,����&��\��Lbdѳ���5��g�D.�b����Z��Q8\8� �%��^x~���-<4a)r,��0���n�s��\���{ﮍ׾ ܏��M�=p�w��O�.�L!sVI\�f���GB��|��ٖR�$RJ�|q
����oj�H�w4��x"q�$�u�� ��u={M��V�0d�Î�~�����-�������T% I�����4�X5&1o�G���y'����|���h��I{����x��a��i}-+Va�ϱ��3Z����c�E����޵N�� �~��4�<Pz���:p�Z3u(Ҥ��` ZV���������Q��uǋ,�zVѫpO�~�u��A�$��[��&r�vZS�/׊���De��2 /"X����x�f��ssV�/��3߰q��\)|v}�L3���1�\`nA�)���k�X-�Ѵ��~���Og�>-c��g�>�P�ǲ�y�)m�XC�+�l.�7��r\��ۛƍ7O=qsK%4��p�ce���3�|��1k�;9~�<�_��ر}��ZX]ZAwϐ�kes���i��9��岁y�X>̍�;0��R�*�<kr]�د��\�$��Q���\�ji$d����*�{�VV�ճ�h�ƓH0c���#��oڶ��s��_0��@��J|�o��������Z)� ��}��b%'���Z���K�36�<}ެ��M���&�W�Sx��~%I�t�z҉�U�C�ർT��:@'-I�o����{ݛ�{&"%���G�w�<������Ő<�`����)z���l]��+�Ҏl�hlm3�r���w���q�*��˃��W�* K�`�Ҏ�d�9�~i��ѓ >. (�Q ����4�����>�����=�^G�ܚ_��K���ډ�������yQ+a�架EǾ��,`�_�O���^�䯯�~��S���.aM�!��}D�m�s�iL��\ǟU���^�����W�2Y�Ύa�A�p4�s��h\r�عs���x=F��X���j��춮,�kqQ��e��"AX�ک�X��"���z
�K'�3�;�S�,?VƗ�{XJ��|H$��w�)����9�ྟ��{��)VPc�z�^o+�H��������<y�~\��7`�K_���n�z���,��:�;��{v� ;9��L�c�T6*&E�6��0DD�^Ğ��18�1�hUT�>�D��n�h} D-X�����,�V������Wׯ��/����d]"�������N�f�j����s��?���R-M��9Ⱥ�%�m���ϋ�㊢#�9�*�ѓ(x��d�&�20�������̔
U&���]`!��M�A1�h�
�40��1@���]yF�I��������gXb�b0�7}g�+2=JISs��]��R�~>5^���Z���AU��5\1y�g�� ۃD|^����>���!�H�W�1� �N�������&��{��zK�0�:��4�����}�K�ӱ���:^�4������snLЉ�?z��[4ѨƠ1������hͽ�C�!0�k��M�A��(Z�X.���D�����K�{х���i�����|x��8f�����r��-jD�t0j�9����o9�V��Z�"��`���E!��gtڌZ�&C��$;�7��?�o�cG?��i<���15��r�܂���糅 �#��������y��'ൗ��y�+,(��y˥P��>�cǎ`���6?sF�����JY�e�E���]��bd]��2mS���?7�|l&�T���60�8���O�lՐL��ח}|Ӻ�_{�?/>)���l���_��O���__�����h ��E�[0C�6N�PU���7�I(�
�%$�"?scRk���k�OO�I����Ŭ�F�z�����SFq0��PŴ8i~%|x��3woA��&�Ο��x�9�#0f������z��0��|w�����W4���h�뢎�Y��c_c��x-����������^s꙾�/�'Ѷ��7�h��S��u@i�:	3^�0z��7>/.��-O'^��u�l\���~�Y���שxAD4�g������¯����y����j�kYd���U"*LS6�m	�4��������+_�J�! mݾjM�f���70gcZ�ˀL��a��D�R��,s[��L���E��S�C:2�D�&���p�F��E��?�S��3�;�|���#LN�au�R���,�M��uCcV=sea?~�\z���K/���d�L�CC�����ӏ���;M&�ӧ�l��W�� J��pk���SN݌�������H��ɔ�>;�³?��<-$�^���o�ƀ�Ց��O���������XL{ߜ$��.��[?�ȣ�_]�S���MA�mb���o��p|�g��6��}���$^�n�II�������k^�צ��k^#�J�1]�
� iܞi�X�n5�83�O������1ĸ����B5�����f�ǥ����6V,g�z~�����_ګ �h�rk#&�?�kq���c/8����8�Ғ��(�f�56�f��JGMwtъ��_~�1K��b|�?���($���h@Ϡu��Jk�b���xZ�wF5�yO���L�֘�p��Ix��ş���1'~/�9���B�h/�I�;���R4;�X�ȑc�D�Q3?c���K,�� 9�Z�e+�:3=�CG�Y��J����NJ����l���禬9��U���>Ԅ{z��u��@�p�$�I�#B����¨�Zu	��o��מ�{�~>���Oca1������Ba�	]��CX7�ŕ%���p�Kw��6WW�)�²��y��s�?�M[6`p��KV��nX��L��S��x���2�+ؾs=6o�enL��!x��E ��XR�Xjay�����sg�9�d�$&�f���}d]��l�=q�0����'����+�|��>���^WfM�L�$M��;�y��k`���I ���X秨�	#q��}!���U���3�N����y	��x~�l{"0�_�_LQ �AZ��Is�A���ύ$�0�ʏc��;p�{D��"0���l��缓�����|~δ�vB^8�@�Q��5�O5�bє4U����Ǡ�p��N�(���د�����S�,�^���F<�,.��F ��J��E��~޽����k���ʇ�+~}ԝ���W/Ȉ���(E|A{����+/`�v��W=�Z�Q'@�'��`N'��}��Sp饗Z�y �fƢ2u���.k��{0�̻r�f���Y�8�n4�~�\�����h��������D����l^U+Ze�s^z6oފ��)+So&�SӇs]��Ew������m�:PWp���عm���_D�Ȃ4-TJ�iu>| C�شi=�&W���d`�9���Ù5�I�����!��+X��еh֚(Uk�[����zt��@?$X��@��u�\��p�������u]w����<����s��m��+_��ώ_Pmf���%-�2P�OU`nL!JM�!�(���#���^�t���;i�w���h<�Ƀ.�k�Iz�" ��/F��ײ�U{�'���K��Cҳy[c�tL��K����T��92���E8K���ʽP"0�@陻 S\Ϥ�Z�@y�7����g	zZ�N��g7��ĸp&S�Ƣ��@?��,?��x$�VY�6�<��)��
��u�?ן�iRV#/8k��%���	��v�t\>bh�УϚ��$8���{���'!��DS~����ջ_l.�����:2����_nQ؁7"����	Ԛ-��)�hf��~4Og����Ӷ���|�b� ^3T���l����+�� �h1�$e����2R��k�4R�n���景�R�o ��1�����\�l!��'Z�V��~]��Ь�Q�T�j0 �``�=�t6�]�v�7KO3�U�M�H��?xa${6��6�bI��}���MU�ZC���Vy�ڸ�UC6���Ʊ��ۺ�������x_'�|j�u7|冣���)!�踈�9�UD��� G`΍C���7����2`"\��>Z���q�߼q)�/��1-11��T��^��İ��(p��fM�A�Y�v��H�ǿ�3���<@�����L�ln�0�!�}����^�흸��g� �	=�j<^0���I��r�v�+}��?�4�cHgz�\���=-蹤��YH\���A���~4f	=~N$��:^8�s���婓�#ˁ4��3z�F��9�υ_��5,]�c��I��[�~|N�{\�{�ҹ��I�u���;<�|��:!���Vl�7B�ͱc���6ȧ����G2�]�ˡ�#�95s�y���i�6uXc�t=�eU$`Z0}沐�h����8h�a���7��Pi5��$Q���3��������YX+����w���R9�Z��^[A2���|�_c����e�*�`�H�w�h������T�(W��M`NP�V�j�J|��5�h����ו�5<"�zx^��+�1XsM�U�&>�ɍc=�u����É�/�"~�40��}�~�K_�YyI�4j�/�%���Aǵ6���
���y�|P|ύB"����d�f���H���W���K�b.�Ȟ)j3s�rC����y���HK��X�L���N���@��351�����*� ��U����X��ӹ���qF[�������9��&�f�Q �g�:'. �q��	�86�EHC����<ާn����M��1q�@����S����S{�ܳ�ߵ��	}���(���ךhn�o�s/�z0�����~�=z�D)y�|��}���$���c+�c?�^��_��-��{S���<.Tx���0���4�&l15�j�7B^9���� ��ulݺմI�����{j��`�W+vl#rc�&��Z[��u��P����ۇ��a"��S�n��k�M�g�A:t��|�Ě�;Af5D�[q-��nU߭�C�h��-X�+���+s�����?�Wظ��+ed�A�%������u֩���UY)���q�I[(g��h5v�T��QJ�g.�\��?hۊPM1��٢@R��)��+�_���\�y{��w'��1�=���w�����r˵33��Yˇ��Q�V�(�}��%�X�¨5�"m����4Gm_ K��מ����򮮜���. �`�c��N����T� ��faf�(��k�bv1�8C�g��D�4N��y�s�Z6�s���̕s'F +�)���3M�;n��r�P�[�]�O���]@�g��(�Ѓ���Zђ��_����Ȩ#P�{Ee86	���iTh��7 ��`���K(�M+����p�����ă�D�	%��� ��B䉬D�g	bx-�)��	�K�W�F=����U�U����ղ�{Te�y�����I�����}����^��xm*
<'T��JҒ�]#$6K�q��'�Z�Z7�VBFM[�̆�2���N$��5�"�5B/t�;ep�����-B������\m�M�k�?JK���2�Y;��@c�����adʶ�Q��p�Ȓ�I"�����N��J.S�?�����=#XYf`;��,}m||s3��>,-6q��1T����@�?��l�j�m|Wƨ�k*U���ǧ�H�E�s�*�G`�}.�f���R���-c0ڗx���O<Y��{�}�_����s�����g"3P��F5�Y#F`^X(�K����PE����/�Q�2�������1���9�c3YKI�dړ�@�) xxFﯭuc��Zƃ�W_���q�9�1hn��:���W1t]�?�g���kkg��Z\s:����'a�k�^X��=�Ƶ:]��m u[��O[�p ~W�>��#F���Ӹ���ki~?w�G��@��1ᨢ��A����^`��%�Ư�5���]��Os�Ůȉ�<�k�H	�G�ȭ5�z�2�qj��0�9�u�C�
���v3��#�=�ɏ�Ԗ�ӛ��ʄR/����?�9_cc��+�t�f�B��b�>�F�����TH�ܴi�YV��p	�kd���<D�hU����.e�o����܁*k�;0'?�9��;E�9S��ȧrȤȦ�x�5���gmE�VF��:�m>�;�Ʈ6q��$J�jTbu-`9�i(NEP�Fh&t��-`����Z!��]|2�����<$�Fo_���}�uC��_^��O����G��w7}����T]�9���XTn�=���e$��O������o��%I�U�j s#�X����B�������6�5@iV�f��T������ɺ�m�(-N��g���[3�	X�{��`����k;qb��s��H;�L�Ls���kκ~����Z������o��7ϐ���AJc׼y�Џ�3��s�1x�V�X0Q�]�6�T��s�xzQ~�����8=�q�Q�wE�{-ү��mOk]	t�M����|{�Y]t&@�P^����:ѿ���h�w����1�f�
sJ�2�=���nO'����Б��$��i�1>1��|��_�[��?�5y���~lܸ�,����Ԭ��U�/���8O�L�m�����K�M���¼�rDü��h.��(0��ڋ'�<,}��������l
�tW��J�w�)��WQ-��7`}�Y��g���9���#S(�X�j�km����9��xx�gΎn!�-ʣo�4J��Pm���9<6��c�������I��r�/�zǝ��\"�w�m07	2�F-��	̹P2�����i�R]dnB�'������$Pn��@�B����b*b&���������bҒ<��fz����:i=bVb�q�C��k
@��yF��ğ՟<DP5O���f��b���S�=ş]��{p��}�<ƛ���'�0F��A��k���/y�_W��9qpSż6�D��^���=x�� K������ڦݨw��5���N��ǧ�����>`K{ħrʼ��4_/�h�i��YT�+��ׄ����-?F����9�{���	:q�DZ<��m�#�/M ��ӹW&&�ۚ9yycz�vV,��3��r�,W�c��s�ְ����G������[Q��	~qڷ���p�A	��|$zO0��s���LIV�K�z�45��}@�<�I�+�����z��ʋh6�ؼy�K-,-����w�^��~��,�Wʨ՚HF���L�	���.X}����,(��r�4*�9�z��;�~�����ߙh��|�C���O
��.��_��������R����&#�dT�2�fB�qM;��#������yh�3A�/$��    IDAT\�\��Is�,��#�.�+`2���̢���}���g�Ҽ�M�m'����9�ků���<��J��H'����ڏ).Lh\�+�5c��3���%:���܃�?Ws�����?�����/Zz�3�->�/:�8a@s䁤��&}��� 2��~�R�.���Xs��j�8G^h�{��ص���9��d���Х����ܶ;WtHx�Fg0���W�"O�nf�E*�/�,LF�	�L�:	E_����y���-x��Td�����op� qa�2��T���C�|��gXLF���F����G���CT�Q�r�upfv>G9��&+e��(n(s��K2
>���4�{�^\y�EH��h5kV$f~f�
��� ���Z��R������T�J��9��������X�*��S�������o'	5>����'�g�B�������w������\IS꣙=�5�/R��I���毐�75��i��Q
�Z ߓ�E�b�I+��2����O -f F���l���N@�kz���6�ר���W���CW�ˬ��Sו`�	��5=��r����8��y�Đ�����S�u=����[�y�	�5/��k.�x��$���^d:T$ ���	.���������Γ7{Bc�zzК��X�i��P���হ�r�G���gH����:���ku҄���� ��Sc����ka/�6D�����`~"���B�������.d6�H2����`~��1,��d`N�@mB��S��M��̼2�0�d`���z5tN��F'������F(��.nnW̆efG5䏣���Z���H6+�d&Y���F>xj�4��-�?w~��עժ�^-�����Tꘚ����zl�Ї������
��t4֫�j'sy۟�.`�*v�ۣk�����׭��m�r ?@��w��s���qR4s�e��+7�Ǉ~���%�4�s���2����)cn��5�?˜(0S!��WB�Զ<'I5��I��a�yyMP�G��31H��x��P�(����3�8@��Ꞓ�= k�_�)V�����8��Č= {�������9��:�����s	��똶���<��i'�<mZr5�9^�ވ^ǹb�`���8��>^@�&��m!3b΢O��P矗��B�A���p<�kq,��`����$~}=�{������C޲>��k�ؔ6xmi�Ap\k��i��s꽁ntO=�h�R)�3�s� ��0��S��~K�Es6E	=)�Jw@VS����#��o����6������h�iQ�&=��4�Z=�j�+3F��6�D��9��S�e^_`Δ��,�'[E�������Ch�ڨ��P@�T3-|ff=}Cضu.�ӊ�D�8����a�bI�Y��(��^sˈJ6���t����uC�m[�7�D姁�����ǖZ#_��W?��?��J���K3�`N�\�L����x�J3*�݃���ߓ�L+�G����Oy¼%]֑��37���h"#P2�R�9�g�q�?�^��у^�ȼ��Bb�bܚN$=��1�i��?��h;	$�/�J�E�9��_��ŀ���|��J����@B�k��X<�(;�[�iGEGn��� ���X
F	|�i<���Ȯ�N����)��~�k�q������,�VA/.p�^�n�]&t��{�N3]W����֚z���4ma����kk�B��h/�L���`�I���
�-�-�K�u�T����BfF�f�u~���mk��!+�P�B�q��NK�2���r��g�S\-�Ϝ��&E���eYSDf�r����[��б.漿���ed�	Q�)4Z��(�^:�3�Mg��i��'ϧ���N۳	���o���L�@�;[�U:|�]}ؾs��`a1�9�����I�L8�r�sZ6(���S��=[6����7���OY#o�!��^������u�=�«�%'��63{�ѭ��ml�Q��r�D�5477�џ����H$Z~&3-���F��ˤ��čB��!q�~���yH�w�krLB�F�OK`$?!7����#Q��+7�	�tt�UԲ����ĵ=������p���o~][߉����m\ ��i����\c1o��I���ω�[�h*R�4�f����AӴ���(-߃#{D����<�Ͷ�����T��uE3�+z��*�&*Q�	�x�Q'aǃ�_�v��;YB�`(&�q�����\�,f�k��ZO]�z��^��#���;��C�.@kJݶ�4*�ۗ�����=��v��_�1��in��xϛ��70^\���b�9�K����uS����^����}}�
��q��y��0k�Z��b�c8Gz� �sT�ف�}�*����Or��ǙIf�Oz������*�0��+��\;����?�nt���"
]y�Y,��019�r���{wb|���9�K���/�g���Bkt݌�YyF:iExZ���z������M��%�%�O�uR4��K�?���������5]���BO(7�r��Ҕf�.�яZ��F^���	rc�	��8�p���eR�����(����I�������&6�KÒH��LIچ4'1V��3Cњ����ך���P�9撠����N��UEL:i�~��{�����'��K�J��F�M�'*��'��i%.�1H c�y�,m]�eeH��k�����b�=�$��+��ޗ�����h��mtÓ0@' %�IK�(v$�6bW�&F3�Yi4҄FfvdI�h� I�$C�&@���=�ޔ�JS�>7�}����Q�bbCE�������o��{���f���J"�t�;9����/0㾜7uiMo�o���c8g���֢d��c���hF� ����UVc�v@�~�H��Ո��b���=�w�5
g��ũ�#W�e�׺��pC�	>j����T��`N7
�� ̑Z�2��^]
���b�2
�P@��q�D�34~����H�`�sԼ�p��h>���j�z-_:X���<x��}}�x$�`т �Br��t\
�����o��/�@���WwR���biQ6oZ/�3�����%���efCu�{��9E-�����h�]�ɧ�����S����O&������,������;����
C����wCe��+"�6�5p�R��d�  ����|Mv-�����_���m��aÀ��{h�8S��=m�
{�^��m2_͌&Gޖ�ZFA�QK�V�	3۰��E��`5� L�I��9��)0XA��L׎�HX �g!�k�i�;�]���~��ƿ���9,@�y	 �ݚ�񻥝��\'^�Z7��鵽Ϝ�D͜�ӳ�� �>�јH<��Aవ�9�����&�ta�D��8^΃]O
>�5&�Y��t�9��
������@0g�����z�}��4�iIV��k����d��a��rL�
��ĳм�\s�	��}����4�م���*��]b]�6�d3{:��)-w:11�����Oղ�my����w�^���sk��I\+�Y0� ��r�tTz��϶�㋲z4��!^@�F���ܢLO�����T�m9rlZ�X������O�^6���\�����ˡ�|�;��
�ml(�����?��.`��[GO���}���G�OE��d*��\cn�`����qv XA�Јif�;��o4#ڱ� �ln ���ZL���ס��`��3:>ü���͞�5pOl4���0�s���J�$Ȁ,qY�f�$j�Ti&��Zaf�~`nS�8f;j^�-�'pX��0X��N0��b�-��g����\h�Q6`�oٹ�`f�@>���)�3�������t��6��9�VP!m��8���W���X� �q�X hi�`flṠ%��9���(L����[jƸ�us�9\{o+�ٵ	4�kj��9a�	wl����N:��ׁ&j{/\�t��j{��1̵�W�#�s.O`� 8���=�nn\]t$S�5�'��sܷ?�{ׂ9�k�qZ�>�7��c`Чfn��DԻG��P���S3�MJ*Q����_�M���M�)�&J�Ƥ�p ��7(�VL��J���J�Q���>_7��8��՛�T|�@_�_�w�"��\�g=��̟y��ٻv�y�����(�0G� �a���#��@���Z����n�8V�J���m[�mf*��g�&���Y]7����麹9������/
0�2�3'�)���eP����^�jDV�_7��^v,�V� �Xf�kZ��	+�����c	6��5p�����B�r�K�W|&˔��±��&��!P������6���V0V�����i.�9�LLm���)�R`�FK͋4�%����$�ZXa�����l�l��ųѺ��Dx��{ϰ���g�<�'5��:C/��$���s��uX�Y��=�¤�1���ѫ�0.]�� 8\on����sZ-�SHR���uЊ������Vc�s���li��PO_��}|渿��1����T3��G b,-�|���cқ�I6ٔ����ʩ'��l���m�����$������R.U̵�zԥ�v��"%��Eg
����z�t�X��C������߳�[�~�7��*�Ч6�ɼ�g��Gݰ>�;�7�`8��A\ p0	�����Dm�� �`r 4:��:߹^�	5aA�g�� ��|pGiE0U�A�G��D�촄n�e�d�܄�h�4m�^�yM��,X��2.�"9N�8�j���VZN��Lu9!"|O;g���d�V���2�!�jw[ᄚ�%;F�h�A.�� �T4����k���p\^�5��u���&]�u_P��`�5���k�H'V��´D�4i��0��P��� ;����\#
t|F^��@������X7E0|�EwF��Zuqa�����A�V�0��<� �x�/�4�vf~A-+P@p/Z��!�H�f+�����7wݱ��\?�]�/޸�����m�=��^��3;���<O(��2I��E�s�M�^&;�o��4	��=�*|��KR�6%��ge�T��n,'Dp�=���J%�����@�_�����������ěW|s�w��Xi�C�:�9R�\�@?���F�v Sp���$���d e���
@�9����g���h��y,�@���j � $���k��P��I+����Q8��/n4nJ2H^Ú���
��A�W����*�	|��r�,�׾[��� �Aaa9��2M܇Z�������x�5S��y]�}�s�qZA�
�f�u���1-+x�G�}2��D[s����~�q����Mz��l�/L_a�'���,X�5�4���ح��ߨU:@}o͈0XZ3��i������֫[�'<'����w�/�/
��v��Xwט�9ʹR3����b��B��`>=7�n�e `����Z�\�9����p���5�V=��X�S{���� �L��kZ��y�����I��;�ƻ*9����V�� �S�T ��TC��d�\�sDZ�E��բ��f��2=� ��A�<� �E<'�(�n ������E�_�&�����36�^�y.`����[���jgf������n	�|Zl ILOf�R���E��)ia�AS���Eq �7��Tu�|�DR1"K]�A ��o�\P��ɜ�FF�I�c����4*���Z���h��e�V�$��)��,H���,8��-�֌l������a�O �`a����BM����<9�
���4��9��k��d5g'�,�0�ZfI��=_A�]�L�5R�`�Z���`��\��m�lqW�B�WFFG]�G�7di;����}6�<�t�S�����0]��a��
�aAΎ��Q+$p>�;#ɭ��cq���9+��gׄ��M�+�Y���D�2�E��@h�&���6�&��Q�@���H$�z�0�O��)��Bfv5�{�7בZ?ڠ�յ�Dw6ЈStܾ�i�`7��	ܣ��� ��KM[��n�>r��HTA`�&)�dZ�ٔ�3QI�k�������.���cq���J�
bGM�=� ����TE� ��=����!�>�fb�m���������
$?0����>���T)7��(q���Z��m�n�E2I� R6(��0�%h���ۮ�:�?����4ߣO��}u;͠!AX��~9���.�(�ڼc���ʬVL��fl��G
�'+(�Z�gKA�j��F�:�I��0Uo9���k2ܛ�c#X[�&�v�>��4[ui�[20Ч1���r��mN��d�����DhC`���u%h)� �=KՊ�2}6�A�Ͷ�qTe�͆K���]�i�h�riQ�	�gbʰ��yE�(0�l*��Ar9�miT]�4:繒�����
��tVu�Hh���,�|IOQ�	�L$@c(��(��;�k�._�	׳���qM�C��Ԭt"��hl7��`:�9�v��t���ӝ��P���
f>����	�;i���Y�7��!n�6\�c�B6y�^��>h�[�P2�I��p��R�"�����)Ų٥���)�1��4Q��	�mߩ��A[�龩��s
����P#�I�7�)�wJ?�` � ���U4��bI���4�l:)�\Z�鎜�y@���+%��Q�ߥ����BaPJŦ96+�Klw�������b��L�㛆����+�N'~�w��ݻ���J#���	�����]�j�@������;� 0�Pc�u��f�yV��&����&���B�e.V���6��ݑQ8������{2H<������\Y���8�܁F��0��3M�s;���L-���"�2��~պ�td��1�գ㲸X���J��O�~�r�5Q��X,I>�
a~R��tZ��z��\Q �p�9`�����a�F��@ d�Y�8_�'��6 \].���j�/� ��Zn���qc����dRiIģ�k?!���v��������
R)�%��i���RY��f5�I�g��~�fGZ#�Rh�1��R��б^\G+�"Ϟ��S��q��0��iJ�O��o=Jz�?�{=,��}�{̘�q=<�U�ǹ�\�����`���Ǻ+����E�[iӃ/��~�>8P��|(-�V���t0��KJWÃC��?��Ux�Ah*��G�|�yw|�N��]��.�.��m�'r� �������<�w|��@Q�$D�G�+=���)�������M�d����/]���D��<��#��$���
���H��ۙ���������H6d���F�0�}?�8��t�����o��S���R#�@	�9*(����C������-s����#�؍k7�D��g��dM	��n%r+L�wW�j�Yˬx�r�}>���g?�������>�A�3�3��2t2$
������L�ɵ"�y�Wx�q���q=�צb��:�>;�� ��i��k��">H�j�!��,��:�TI�(̜���1�/�U���K
�8c��
�� u-�1:�����T����☙2A�\�ׂ&>p�h.r��ka��Z;����l�d����+.�^σ���7 3�%)�����ԛ5���t�� ylЮ��Ľ�v1(�r��a+hY`90�6Fz�%c.��B��@Mj�Ҧ����ۿ��A�� k�+��g�+�#�s,j��=�9w��@84c�!�\�����ӸˋU�� ��U��u���.��	�m��D��ѧ���y�<N}��MZ������4J�wO�ǰ�,��m]K�Z�� ơֳ$~OH,A4���R��s9I'�~MA����%�t`.X��c:6� �TA�*��Ĝ��7<�?9�����a��S�g6���_��^~\i	f�|��������|�/Wk�7�:�uëx�@��C0���r����DM�޾�^�����Ap���ڃ�z����o�4hd\\���%�G-��Ԏ?,Ą5Y2h�s�9�W+d����D�~VKa+��Lܦ��ߵ�-Y��m��c�d�ȳ���`���!���k�^��+���zQ�3    IDAT��i�ڝ�=�t�1l��L�&�l_`}d�-��v��kSh�F_�.�o mh��C�3M�p�T���d,���'�R�ۓ������U2;�(=�����%<���j�h��D6|��]��ҷ2zo���Lڷ@��h�PhU��PQ�&Z�$�C��+]�@8�Έk� -;�6h@(�F�}�8�����L8��^ÞK����{m7����E�	Ч�U�Z���4oX�v��)##�s�}�wV�C-ug��9�q��:Ev�X��
�o��s�R�:i{�<�{�{0�����V-!)ob�kn�S� ��J���+�D[F��򹛮��^��i�fЇ�LLA(NK��#�\���˹Bb���s��t*������^՛~k�q�x���ߝ(�|�{��ܞ׮i��k2��Ih�X4e0H��s2B�޹���A%<����8/�ZFCD�����hᆨ��<2"jFa�a�i���,��-3#3}��	k���-#���{-W�%�a!�c�{��,(d4����{����5��.'�� ������hD�#�<�W������Y������s�E��㆙S0[\�J2��b��)5�RE:��izRacR.Շ�m��[[
ٜ��(\�L&�qZLD��I&�R*/H"偸�t~�hG�٤\p��2�0��:2�Z��5Ig`!�]��RiA���x�3�1�������2	�הZ6���(I�W|�8�v]	��]A���k5�Pm�H �ފc�I+X�/f�PF��N���.>���B}���Vy�风k�_�����jC��8|Hc ިm�c�Ӿ�(OJ��Q�F�v�3.u4%�&u'9���^m������.F��Z�s�����8����Ax>'�:g,鄖d2��kO!/ٔ��PL>{�e2:��ɑ���Ei6�J˱�����`�0�	.طɄ�ߴy��U��=Dp]�1�8��qpz�������k{/m����[0W�ӛٹ)����j��n6�(A5�0Ҭ�F�j5��ZХV�{�5�(�����6�#{n����\�gاn��@3�R�=�����
�y7�?��]�,��ja5��ظnz}_L#�LkR�#���hL�f悙 �(��3�&�`5j�um��j9�#2�_�;�S���bM��
z��͎,-Ue~�(}�r�9��W_�g�}NY,,T4(.�[W�e��-X�u?|Bʕ�T*e�>YG��­$�h���t2+�FS1�;ϑ/|�F���o�x�����ܒH'�&�6+E)UʒLd4�c�i��k��Pu��[ڳ4�����Y��� g���Bq��_�[h��Į-���,�o��@�� -8V`EV��a�'(�c��ٻǺ��^� fV�価�dk��mZw��<�KB_�/�Zoi}��G�%��TU���ϖ�nV� ��Z�?��Y��<β��8�'��ш����Sa�� �u���wg��\!�ǁ�)����z>�`Z��f�DvRB��"��	)dc�j &�]{��]ݣ`��I(B�/"3sY\lK*���ْ��U��j�� C�ӒD\&6l�qlU��+����8����܆]��έo�{�|�5�b�\7����l���ܨ���̃@Ln:n~�:����m	�~Gf0o��1G�%>,|P �x�:�@��/�����,��{���@AK6�H=��Z8&��8�~^n���)���XA���V�cU���h�l>����}��Q5KBkW���=�.���M[�nV@�W��� �t&K�h�����֮]/^x���λ����,Ve~�����FD��rZ�L�9,�qBC�Ғs�=W6o��ҭ�oޒL&��+�R���o&���^Y�~D���.]�MO� �Z�%��ٿ��y�^�D�pAu��(bnqMh�(_��=x.6��;;Ҫb�\֏l�����P+O�u9�Hw������hvj�q���:r+}�xh���m��ww��q��L���,Q1����sǇ8�,��V����A C���i�&ٶm�4jH�����?vt��9����=<�V��bM�5��M�p>r̃�c��s�X1�
 :~�^x��B��H�4~
S
�'$�O0O  T��!h .�T"��i����O_"[7IL��j��"�X$&ӳ)������\Y�K�KG��G.�A���7�����h�"����V̟mj�m��í�;%��10�׾oo�����ٹ�I��t��'�G�!��!R#�tN�!�`s�i���52?�@� 6̬cK4�2>�	����:>�l�D>w�FX��<[P����X��s]� x/065?F"��B�#3�s�z9룄���2��P$�ש��ʶ ��eM]K��bؔJ�$���52�jHj�j�Ϯ�/� "1�ԲE���@w�v���)W���r;�hG���뭦�DD+���X)�/�W�W�n-"�&�L�V֊����Ǝģ"�tT
��<���z��N������bS��^��ҼjKҁ[�iU�Ȱ�̧��75F @��bmwjs����3�D���vK_V����rˠ\E����+�?��F��;t��5 צ �@�S�`�,1&�\U��X)�A0�v��zb��8��ޏt������tSC���M/���_`=`5R�ZQ|Ær�Juq�i��@m�F��ZZTzi4X�1���)��of6p}]=���68>��`o� J�;���0�<i�^̡��$�>��=&1�er�I�uԐO}�"�v�����1	�,Q��[������C2=_���Es�!�E�?�c�Vuݚ�__�&������V̟y����z�-�����#���������<0U���p	X�d���aa���� ��s��ڀ��`l.�*Z���8F�9L4���d@V�	��
+��}��y�ף���ɛ�q6u S�>v����ǹ��I`��FFIf�����@S���d�8��hQ���8�c���ϔF\�o`����fU�6z}iQ����}����3垻�R�=y�ZL��;��g�yx~�-�����(���KoO��}�=�o�i����$����H-˥SR.-H:���O=E�3�ym߾]��u
�ӿ��!�F:.������e͚Q�['�?�G2�A�(̴K�%��ⱔ�` M������K/�\a��C�"���c�=��8����Y�&h�K��7K/J�q*t)a@[4�s�Q����J�0��+Ǜ��6��/"�Z��2���	Ρ���b�x���z�s��Eg��h�f�r
 ���`��c�(�q�آ�%:�Pk	2'��7nT�h!�CDjժ����Oa��F�fP�2R�T�� �ŹN�r7�.�{����h�F��[*&.7�ef���@��+z|:zJJ���℠*���t���3�`����[Q>�ɋ��3֩fwi���#Я%�%����P�`��t�����u��!c���ۖ��aju�~�Ċ���O�{�m���f�'ai�s��Fi��%U�i��꽏l3ؔ*��%^/l.��U��p���p� �@n5�0�[���
0��쳆A��d���ĸ#�ٺ�
 �Z�|�.���Z�Y��k�)����`����c(��`������N� ��ݻW�;'�p��!����)d��Bo��-F���B���T؊J!�����B
��|��_��k�(��3V*%���	gq��'������ʍ7�,'�8,��w���H���H4)}�5��f�$ب/��������1�w߽�� m>H��ݤAvU�f�����w�#�^ �֌�|�R9y���dp`%z|?�y5�v�0A:!�ګ������i����2�+H��C8طo�j�8�+,�Ƹ7���o��e��*p��z��@r%�gNa�ҹ5SP����+��16�V0���{��p��,��1���q�1s�:��u���u��@s�#���FU�%!D�#�>���Ӭ��5��jͥK�x*��2ʼ"�F��p�=����:q�s�[�D�M�@�
,R�8�� �؛�d"����h�U3�� �x<-�H\rل$�e��s�N����HuWM��ؐ�bMb�K5���%BH�7�/�"u*�щ'�_�H��?į��?~��o�y����.n��=�M+1���7v(�\���&��ЭFh7��0йMG?�+�j�x��yJ��<��{��c��&���A3�������-dZ?�>Â���V@�`N��-��������Mi>Ż
>%���Z@h�c`P�Q� r�eAk3��/� ��>����o��0#�W�4��#ɴ���7�/�DRt��f����4���_*_t���˟����O}NQ�!"dc�	#�ں���2>�V>r�e��x�r�-��K�H�S�����G�fP�.�ZEn��z�/�)w��my���dq���T�yF�;��N%Q3*c��r�eJ,�L��D��c�Joϐ�9��مY�����c:��^Pa礓N
:b]����qnK����j�`������u��hv��r�Z&V8U�p���{�������?
�#�"y�Z�8^Zy���}D:֘����2���{�w����
�����֢5�{�3�ȵ��,�U(M#�=���êdy�1�;�hq��W��
�ܗpqLn��*jn|] W:O�tZp/��О���\�����b�뢒��%��#�tJj����u�E۸oLұ��W���l�k�ޮ`j�93{�֖�IX��4`z�$�F; s��x ��|m���o�Zq��>į�{���~����_���{{�*�9m�������9%j��O�	���5��:`�҂�h7�մ���k� b������%D��-ྟ@q�����"X��-�[��
,4#Rs�fD;V�C�hr �d�xfO_��'��l|Mڈ��Lv��Z&Ƃ�������g��I�򩱄cZ��Cj��5r��!=�r��9z�|����W|Db�����|M�ygBʥ�Z6m� c#��7��v��wp������j�Za)x��45"q�����Ų�kF���?w�߭^=*O<���291��r���~�ɷ��FM�l?�4�����'�z1�j\�|c� �x�R�JuI���ia���l�J�>��3%�ye	ZjmԼ�`�8�O�	>0��u>o�2�8�&r�t������B��`]s���Yz�'�rq�iL�-x�|��碶ɽ�c(�Z0��N���@�`�����}t5��:^yh�Z@`9�W�K�+���ϗ��E��}�u\�ZQ���jp���d!$�?�UA�M��c����v-6��b�
q>r't��N!�Z(�T0I������b�#�HG\Y��3r�Md���H<Z�OX%7|�R���jȇ�S��]���)�fze�ޖ驢T�&�D�m
֐7���u�K޽i��/��Df>�8����`~�~��w߻�O��� �p��n�̹8���@��O�/��i����4Ec��@P\N+�f�������,y��3�[���.G�'5{+�,���i�8��y�eh�\2v0z0�ra*�[�l6?P�	��9�4��pǧ�9F�������I?)5�:�u9נ"�E�WTz�
�:33sj������Ǯ�\��G�\����$S�25]TF�����ԓO����믿����~�N�'�zR�z�m�(�k�ٔ+Z�-i����^���k������>����l�G��K�% Z�椧Sr�Gv��kd�5�ԓOʺ�էX*ִrL�X���I��-�5�����WW�)����M����7�x�I曖$�ڼ/ܮ����	��V&�r5�M	��WS�A��	>����5(X��i�ΐ�ޫ-�p�3Yc��d��+0��������Ɛ��v�I/0�'���AU3{C�K�Z�4V�m��O�H�7PE]G q�j�c��O� B�V�w�ېϓ�t�)<PP��ܞ��P�"��{͗�:�B��Vfx��S���:|�VB2iD�/ʦ���˿�����RH1C �c��)IĳҊ$djr��y���$�k����}bӺu7F-�?L߭8��q�c�~������b� 0�)����^}iK_��`M0�Ʋ`�clt��D-�/�a�"G�� ��ۂ�"���IZ�L#|.�f��V�&(��ˁ%��`N�޺�L�/�iF��~f�)có�2���=��{�90����1/Xq��L	�lb�e>�� �{jh�33�jhX������}
��C2<4"O?��j�3���g��9|H��>����;Uڴ�F�}Z��
����O~��24<��>�=���ѣǤZw>[~��z]��gd�	��k��z��-�HB*��H2�s~O�B�u*�%I���O^)��z���g�m�ޢAn�L�D$%�fK�ԎOjT{"��JDU�|�I�.��b�6�p�nq�͒���e��x���,|���h	U�p_�@�����q
��,a��!�[Z׿;ݼvZw,ݱ��
����ܾ���/x-�q��@�|ǻ$h��8U��I4[i5��A;����ӝZ�V��Plㆣ���lo�^ ��0��ݧsc�v�SޙL;��&���Ս����3�#��+.h�H>ݫ{%�IK�ӔXҹ��Zv��TR$�nȺ5�җ��$Z�Ҫ�9Ut��G}{��L�
h��\9]��+z3{6�~q���������y��I��͇��~�w��H�i�0�9'��i�ϜY���,E0��A-�).�`�­��= �k�w7��Sr��`D��K����3[@&�c��C��/�a��X͞m��|��JZ*��^�V�s`{xnp>696'L��!O���z��&"V��AL��B&���v&u\�V�)R3��B�;��Xa���Vw�W_w���U�FUz뭷����r�ȶ�O�v�.����ƛ�舔Q��Q�	/�Vw�mL���/K�ݒJeI��e�ʧ&g�Vs�����;��%�~�ٲ���t}'��宻��`�X<��^ov�ZC���������ϥ�ƛ���ބ��u������憎<��S!`zvF��z����Z�Z�b��ݪ��W�q�a2jj�XG2k
������r�@�~���c��c]	���>s���6���q�3-��<�L)彩���aZ��]�E�s��-�������h������Q(��ɸ�6�3����%�XuI�9������x^�^YעF*P�F6��p{BT����{!ϜZ�D��u�Ѹ�9y�0ǋ�4����/�^oI:�su2ii�jf�t�vTⱌdI&"�JTed8.�����/��70�����LIr��2qlF�p=5\��s]�HM���ۛ������O-o�0���`~�X'w߃���y�w�X��0��&+�1m��숰�WZ7����)X0��1:�hA�� �aCX�qy�݀��Ƶ`N@��F��`�wj
��0�¹d�����4s;^
,�����A�?���
��� �Q{�Fq&�0�s}0g��`�`J\kjm�j-0��wNm����{GT��Ĥ
��C.^;��e������lF��/�yN���rٺy��������1����� �Ə<q����Ž�ޭ���~I�Ն�t}���drrZ�NLJ��l�u�C�ǹ�Y�NC>z�%r�I�un^|�E�񣏫��D�Y@���U��i^(�����?'�lT�������G����Lf%�푉�)�`5-v�h�����R_9�Z�o���]f��D�Ysixa���M˒�L�GTLă�E�-4sҸ��C����4�<�������k1�k`�oaJ0�V�-
s\��pm��-�Y�
4��A�S�����A�?y<�/�%ª0?61�@��G�饗ʪ���^ ��a�!�iJZ���㉔�t��	�]!��K����v�T,�?)W�%����h���A ��[ �g3Z$)���{���ӲjpL�q�h�,����|��2>���N��� ��Q)�[r�Ȭ�����RG=,��;�	֥�&�V��󏌻    IDAT'l���H��#��g^Q0�����������ϼ���T�JJ_�/��+�i.��Z'��A�l��ԉt%���]�c:��,(�kC۷��I��m9"x�o�۩�bl�1�a5{.5���I#���{_	Ι�\�nF՜[N�̐�$1�gޗ��}vl"
)��8`&s%���3V��؜unvM�����V� (X�	M�:;.��1#�Ly�}=�235'C����7�W�]�4/�|^�����N���|���|6-�S:&D?��H�e{��PмX�1���Ɉ���e��w�SN�գk��<��O���ح�ӄz��Q�I���E1���'�Г�_أ~��Ւ��8�I�GP��fB+�v��~�գ#�s�y�������H"Q�$%��j+����g�̊a����O*��~�fP0�>]�V��E���m�9� f�]�{f6���c�:�A̟�
ʊ��P)\Z����h>W�g�A�6�����xV㧠�h�e�@,�s�~a��
���yA:�щc2_,��
јZ�FW�rB�)s�G�^��vlԽi���G�"
)��\� � 
~m��&tl>\*�r�Z�M��&�+��_IC�ۥ�@ ��f�G��eҾN�|�$��I6Ֆk�#�uK�$�z��H8CzZS����a�/.��|Y�Z/�g��*h�ДH�:�fl�_m��w����
���bg��o|�ϟ���M�O��ړ�`���w�Ȃ�2U��r��=!b�0���h^Dz��*���	�dPV_�������F6���Sٕʝ_� j�����Gf@F�k�(wH�AT?��,#"S�s�:`qQ�a͜L
�a]X���h��lk���h��s�}�aAG��S�p��Ҝ��bMٲe�lܸY��wiz�a�_�zD��$���4�}�������7խ���S3�z]�c��6M��������d�u233%������q�R�E��Wޑt�O�g� C@��$ӓ���gzT+�[�	U�b���99��d����7٩K���X��v�a���?�'�T����<��*�~���(Ͻ�vK�p�+�����̜�Rie�p;<��Z��|���h-T67���8��¯Z��ڋ�W��=�������?4s�aP��i�.in����!
�tk	���@2-�4�U�pp_��x������/���|I�`yD ���վ��b��@�(��0�I�Ѡc��8Ų{`�f/��g���Ju��c�t�L��
g�zh�y�9r>'|��r��쩌�hR�\UHSC�:"��7����qL�%���K�m�kI���-�y�������\��̜�di�C��q�F6��������t򖾿\A(�@�jE5�S��[o��W_x������sfe��W��\�H����42j��P��@�M��	 ��H{җ���lA��&�����L��e-c������6c%|��������N�Ei���h.�Ȥ ��q���A�HFLfI�@��*�����{��m�};�8A�gp��z���vD���%j���]�hL#�4��(����9唓5�|r��:m=�P�B�
��vx�)/�BFT�)ڐ����{ߕ������A��.��|]2�����?8 �FDKq"%�X��H{I
=Y��/}Y��RF���TaNG×�RYҩ��-t�V�)��3���٧u_�گ��F�?�����U�k���#��|Q�� ��J �#�
�$-PQ8���ч�lky��V���zQ��F��Z��Y��[�/L��x��,����/�зO�ڦ���.\�����Q�Zy�o+4s�-?��s�\� s�#Z��o!.�׹y�����4����y�j�� V���k���4Љ�w�C<����k�5�����K��A�� j��ß/.�� 곧�W!�� �jE�G̣��\���r�E��Ugp�P
� �Ç&%S���sM��n
K��j��zgh��?uK�E"���	����ZQ0����]����W^��vǙ����w����Q?&}7.j�۝
Dƅ���D�$_�ڕ���A�Tf���Q+�S3�9�
e���-��Xˠ�ħc�k,vVs��p�_�__�G�[Q+l>�g�),�(�t�����L�1�4�[!�jMԴ8��s��[�i���n$h��:����p$�Hv�/U��Ie>>��V���:�ed~aVN<q��x�5�ҋo�[o�&�}���N)�S�$�K�>��jԚ�n���o@5�Ry^5�d�"�f|�����29Y�.�ެ�@Ӊ��&�ޞ��w�6y���z�g��'�&K5�Tk֤V���ǖ�n엽{ߑ��#�ׯ���ќ�K.�DN8�D��?�)��%['��3���ejjZ���x�V�X�E]���>�\��rkA-�V�FH�ʰ�F�#�3�7�V�"|44i"�V�� l����%=BH�����s���/i��*���}��������;+��7
1v�^a!���`~��a�D �7ku9��3e�	�0����8Ar�w�Y☞ب;a���J���s ���4s�*��~��U�@_�S�(�X��¼Zdp�LU�P71;M�a-h��X\�i��/���O�O\�M���a&�A�u9rhF��4h�R�L<3��x���)�,Z�??���߉D"��ԇ���`���[�~������s�LN�>��3���&pDĔ$��Ң�&̠,A�-K  ���y����|Vj>X�va�E(�9�P�$<0��Fa�.nLZ�idp��5SsS��q����G�<� s^S�f�ca�3�{�ͳ64�۬�hL��&�oQ�"%����Ӄ9>;��E��:eZ/��lݺUr�g�Ak6�S��P������u�5����uk�ʑ�����B�W�\�,t.s�gє�*1/$�	˙g�&�|ZN>�9��S�?����'^�X<!�B\bh�ډK�X���)9������|\j�������{�8xL��0延�-Ō|�>Y,�k,���}FV��Үw��{r�e����])�n�O^|�%^-�՚��=�o�~���m���T� fw
EaZ��� �#��8��HX?]�N4�º`���AQKW�q��=g�-7<�c��j�d��E��Pn�#(3��-i��q�3c ק����=j�}@��R��`�V���z��|ʉ.�ϻ�

3����� �նc�*�@�ʇ���}��ۨ��g�qAx�9���(���(���4��y�P,j@���g�j����$Rq�q_�OȤi.ʶS��M7\,�Z���tђ�̏�MV��af��4_ֵ�c��R0/R�߼~�˽���)�;Ag%��7�����~s���mI�f�_�{��w.���W»��uݴQ��$Ct!3���׿����]U9g·�L~��@@�˦�؞��?Mfc��ᙺ��=�ޗ�z�ka��wi���l���$rְ'���ͱ \xoe��{�aڨs+Y�-�65yj<���Xk)�y�fv2]��	�d�(V�o߻r�YgiT\�ГS ���M���*��Q���W_�O}��j�G�%���}����+�K����A���k��

���МW������H�\x�(!��Uy�7t�a�H&�S}�������ԓ7Io_Av��]�x�����PZ��[X$�"�[uG�K���Ko��z��S��ܧmS�,�w?/�~D#}�cD~9:��h�D0_ S��a� B�J����)�G3;����3��� ��`�D\
�/�!��fv
��}�����PP��A�(B}�B?��`�ό��`>P�{����>SK�k�
��c���y�|o�p���Ƴ"xfv��a2�-.ɉ'�(�o;�ĩۧ�[3;�i��#�b�h-���S��`l�����k8 >vZ6��`�5T���am1��VlI�Ы� ���[.�U��.�ߑ!���BK6��/���$����!H�0o���yiE���djfAj��q��{��w`��&۴v즡���ĳڽV̟{����r�mG&fN�C3���wluG3;%YC0�a/�+ �L��2�^s$�GL_|X��u�y,� �oܘ���� �f>�������Dn�1�xJ�xP�axsZ�e��h&�xif�g5�z��L-�����h� Y���s�R�#s  �54^;l���������^�JYk�� ܱ���HgP� "'lޢ&lh��?���y�O�M7ݨu�{0����񏟕ǟxZKÞ{�6Y�n\�I��D^~�����ig�&;v����z�����#����.�ޝ�ZEs"r���b�&?��n��r�g>)##�r�e�\!"��������t"�8b���-��\;1��f}I�n�"W~��j�%�Lȃݯž�~[8$�����J�	S����%����R�H[��
� �X��4��f�ŷ�~[�ܰv6ԟo@�A��	Ҡ��{�T@g!;+��>bܺ�,]Q�kԤO�9��* ��8�<l�b�U���&��fǇ�S��X#p��S|�9|���0��+j �R��=
�<k��Kh�8V���q{�9@�nT]a��U�U����l����ڙ�і�k�c�8�A��
V�~v�Kac)��`��|<�D!(�3�F��hܥ䑩�D�J&.��R��_��+TS0G������#�J�(�/U}Iנ{Z7�>s<M*y~��57G����J�gE���g����7�{˱�����i4;̋4���8����IS.�Uc�c�`�F0C�i�����hv^�`II���4p%vlj���Z{��L	Ұ���qY��憙�Z�Do�n$�N�3�nR�z{0���9����eDޚa-�oZC�y�`��.�銕�qZ��V�w�W�17���hm�;ǉhv�@ɘ�X�7�|C5fh����n�]��hD��7�[+�X[����ʮ���<�_n��&����d��zzz��;�7��+W^y���y�d2�BE�}�5�w�����^�Q9���}�6y��W䍷����C�$��H�P�|�ӟ�#�'��o����䧮����lظV��; ��yI}�Yi6��J��7����TZr-H�"g�y�\t�Nu�K�jf_(��+_���my��gephT;\�o�\-�1\�y��B�x�+�k��fK�V ���fY=�B�;�EK��XO�#�b(0D��`nQ����y�;5o��X�cA�Q�Lj��WZH�D�M�2�@�7ָ����|v����{��x��Q���S0_,�U��c.ѸׂR������ȵ�k�Yvj��HE]��z���| N�W~�=�C�ȋ ���S0	xV��`��P\< Zu'����W�&�pA�GeO��|A{��feU_R����Z4*��浖H&�'����#���I� ���5�}�֛'mZ����ȓ+	��{�(���G/}�;���7��*k����50�-̩�Y����i�0�B d0w��Lоǲ �CD�*�D\
KXy���m5c
-J��P�/�j��왉�u�1(��f�0aX&a5۰�\�hNF/�޼.}�4�Sˆ�����ȴq�j >	�讅�������0�8q.���~�q(�@�F�L����״c"�f[0x!j@
`�n""9�c+"�q��Jw���E�#��{ �ڢ����>0M�Y|}����D����`��ڮ�����r��1������_/cc�2�j@x�������ޑ�*�0���>9�����Iy챟���*���iW����òo�AY����1�Ɯ��w-[[uY`�_r��{���N795!���MA����y����$S9eЈ�f��.����y�`� gXh�z�w��!�\���s0&S�������Խ�F>s
d����ay���-�xV���j�Z��g�+��(�N���t�}��)L�8+pӝ`�����|�� B*�M��E�87��� ���V��4�mO�hs����x��3ǵ�c�aVW�J)��s��P��������%�; �qs�|�|%���S���/���DJz
}�9�Z�4(�' ���AI�[2����7}\�W#���ѝ�Ee~vI�>&�G7(���1�Wm��B	K�:+��y�sd���]���+9��{���wݽ��f�#�NBr=�җw�NhV�꼦׭�d�gH�4bq��z���A�V����u��Y-�n4����3ZM4�-d v#s���,CTm��2/z 9{Fg	�ٰYy�J�~�q�Z�E����UH�`L��r^�@� Ƞ��1-PMp��x��"�@��$K�,��a�esL %wa� q���j�N��f�td�������3����N�����@v�UW��w�� x���CX*�椷7������>�Ad7�|��[���1��;��)��z^���<��BY^�u�B���+�^G������]y��ef���������R�-e�`W7�p�lٴAs�z�	-�9����3���0�LV2�v�*����X�`��C�����Ͳ�ƋgQ�k����A/y��H[��H{a0��`����EAN�\S��
��<a0�=	�>)��V��%��(���(�P�=�l��ST��w;?�;ܨ��N^c�	
!������j��s�"D�u?5�*X�8�T��k�#�^�kY[�K��@X.G��4sh͎/t�9^���фS��C �v.�Fk�S�����׻��{\��7/-iI�Pp�ju-ȄB1=��\��iC�ģ�h��ݎj���|U����Ukdz�,���{���f_�m�c��kV��kצv�$x~�`~����=���ϊ���H$%�B�2(���5s�9ӹ������@���f-fB6�@Ԧn�P��3հ-�{�fn�Z2f-�7;�V���($��@3�+غI�??,h�lbj3�1�1Ҫ��k�6�����������֜Δ���I���o�ߑa�\H�m �fH1�x���� �H?�y��/d��9ͺL��1�Aeٰ}Σr��gjd����;��։k
�:�#��ɳ�����A�@�ޡ�B�ꩧ��~��4��t�)�ɋ/�,�g!���$���і����N��UW\.�n?Sڭ����'���{Jff˒N�5r�j�e���B���k��6� �[o�U����9� �l�z���xvG5o0@�S�w�⚯�M Ǻ ����� ���B��y�v�Ck��eE
�(�-�P��Bu�`Ia�����ߗ}� j>��e
�t�Y�
�vNx.�3��`a��0D0?zdB��*Œ�����q��k�w:�n�����ZS���ܬs%z7��Q����9�L�Q	ˢ���&*�Y0����C�r`ޭr�#�
t%]1'�X��p/�v�6�:�|�W!���BS�|���N�d�`p�iZq�.{��1�[�H��r��ک�S��y$ڮ��_ׯ���`Wr<+
����o>����_�I6�H:�����]0g0�	2�q�A!��@7�1�����MAp@�M�2	�����61�cMn=���h�6�~�����N����ܢD-s�L	C3�`�n5)nd�%�x��9}j~�	�2*;z?�]��J��}>k��ߕu��q��a��X?�a� Pa!Ռfb�*js�\֨Dc�lQy��ɖ-�������.�Pj��j�����h����B@�,/ƑJťTv��y;w�������RiI~p�=*T�<��5���n��s~���t����]"�#/��G�GV��b]r�~�ĒȄ9�'��C�Hm��f0^ �B|�[�R�7Z�b.�Y���X�՚
�`r$��E�,���c�ʰ9�:�X7�J�|�R�����Ej�o��y7LäQ�l����(���M4;��=��Z���|j&}�k^�96��ढ़����l��	j�?���༨��A�#U>s��hvU �Ng��ְl��Y��b�k������{<�\b s�%��-ϡF���c�~n�|	���]�U��AO���q��    IDAT��X�;юZ˲�^5�Ǡ�w�O���Η��m2�9��4�R�!��?$�}�R�Ԝf�B�gg=��k�Q�yF�2����o���{�H��9g%��p��N������?~�س�f�I ̓0&`v��Y���Ծ�q@����x]շݬ�,��p����ڐ����Mu<�w�~��`F���E9Wj�a�%���e;Tt���,�T�=p]�9~#��}��q*�6��hvk�\N��wdd,��B-�j1dp8��ӜI��c��@�9�rt�&���-�I�9��폕�WLN?�dM�:��mr�ke׮�*�_�Q��R��5��d��/�|]�
�@Y+K*����r��ay����Wߕ���l۶M���ި��Ȑ���-��)�*�J/iJ���TJsr�5Wʚ�q-��l�,՚�K�K�ф�)
�0A���<$/����0ѷ�4�����!�-N�8�������6�����v��k�4��^�"CV��1�7
͸��KK۾OJ�
�^�%8�N	�d0�F�����m�[�%AYi�D�}�{Q@��+��pH�1�6�_x.ߏ�C~L�.��J�Px�9x����I�̫�E]�s�=K�1���j�PL��N)A�8��KύG\L��{�\�[�9-X*���7���U���� X:����^�a� Q9.�r�"՚kZ�N�u��=�W���M�>��4�!�<�l���+��$�Q�A;�I$�`^)���!m/�P�`N:q�C0���%�
=pr�o�F"� ��\���`�����޿}��g��̫����8�3L��׺v��", q|�g��%`à%�.�����*��qL��pc+�ht�eN��w��2*�a�'���8f�d�0�[-]��L�7�܎���cͭ��c�%Q�����i30�y��g= ˚��^8���>,ʵR-�hJTFZ͚dsI9��3$���駝"k֮����8�	i��8������W�x�1�H�oέ�5ex�G֬U���'�����Z/���n�Z�$W^u���ɳϾ.��_���E��U����ʏʎ�/ZN���ߺ��Ӓ�D�m�dSҮ5�U+����
�`��FK+ǝx�I:����v���#�t���#.���_  ��[������~��s�g���� 
�������c�Q����-͐�@g�(X@�9�2d��u�g��>[�Cm�4	0w��̓����[!�^��$-���=����˂�?���J�� 8�9:����c.��#j��#����}�(2��P�U-W1�BO�B2����M/�q���R�̓��πy��8�;��� ���_���>�9��؂�?P��k���S񺜿�d��cg"�GbA�s\]F����y6�/�NLf�
���4s�F��}wݺ�_����\��p����N�[w~���~�����D2'�\^r)4t �8s��v�Q�T��B�!6��@M��L��U��>s������y�y����IX��[��S��w���ğJ -�9��7#��Ul��=NP��)���8������>�eJ(��T 0�������&�y.���x�A�o<#5;��;�w��ݦRǙ9���\,��nH:�3N?Mr����^-�3��#_����ʫr��QIg�6�����R�6%-H*���ds1��P[=-g�y�<����G��$�j��M���|�q�6��oK>�*n.r�o�LR.��<i5P���Z�����,�7eq�"�dJf�g%�H�k���n�f�#��^m0ƎgG�:�8"�׭[�.h����S�:{�㹰7 �ЮYP��sM�=���>�< sg�� ]�>#�>��˵�h�%G��	��z���
��k��Ψ	���&�v�Z���R#�V7ޏB)�>�ٺ��|��A����kt��!����مy-�y��e��#h���i�� ��(a��#WP�1#|�0����)j���il�uq�	C�Ν��������G�v�\re��q�0+ߓ�̌D:%������d�UoI!��d�.���N����%�n�f���њ`�N�J$���y�&K��V|��[�!}��#kO\��ù|(_+�������?=��[��TG�+�%�%�rfGJ��i
x��5��GG�Է����Nsh����nNQY��nLt�҆#��H0(�i� ������@jR�w�Y���2@���&��6�@	}��qz_7%w\�ҿ���A5<-�颣�_��h�̔���2�� �`@�O�L���́�=a�Z(��F�b� ��̈k��0a��=@c�v����z��"��u����-��'+�LByx�|����/�P���G��^|E�ٻW���]L�ќT*�e�h-��PVn��Z�U���u9�ΔT���?��h�&���o�!Y(!�,��aQ+~i�,�4��+��ALz�4��fSل�K�R�r��̓��L��Z>�F!�������mMu�a��p
�]����_��%�{`����|g�#S׮Y� � ?�� O0'`[�e �59S0�w����Nk��/��ˁ8���0��4G �#�I+,[�8	����c������|Z�(lZa��׺���/��MN�h0�-���~��(-P`�A��<�����3;�8� ��;���� �=�5���  ��
ت�;L���
��X׺֖�bU�VxV��9�9�҆r��7���T�![��ȍ��T�	m#�N[���sEU[�w�I�
K���ՙ��MM� ��������n<a�/�D��P"�J�s=z�4�������{޸�َI
��
Y�LQ0�j�4ܒЗ�V�L�q�?z���Q1*AN � ��G��9X�ݬ{g�?p�� lg��_���1H�M�D���[��oV�ϐ����� �
�}ое���j���".Qtl�N,*-_W��I�o���|]ՎK=��DD�.lD:��QS&3���5�2��9�g��s�~ن� (�ӯ��`|��c `6 lD�p�~p��X �6PYr�T���'<�D��AK�l�-���q^(�d����4eb�LM֊d(��~�:�Y,/j-l\>k�+KJq��}���"8:1�=�'�fU�@�O.�����ʼ�@��ޢx
͐ʃvB��	�> �Y^,I*��gbLj��[����55N5c���_*-����%���;o��t=D�s������.Z�����cα��GW�� w�/ޱ����I'*�zs6;&���j�6�1�y���id����X�#( P��;�xZ~0n+����(�b-֪e-Ra�'��=�b'�S@ #s�؄�{��;vh�%hB#���N�������t��:�(�hNBj�Ρ�LS:�\�j!Q2��Kg:���
m> �<̌@O�9A=�������V�k���|��֩l*#�}=��Te��Ur�uJ&��ե/
�c_�dv�"SS2�j���U�<�u��7�s�躴��Hv�8a˚/�%��0�'��*c�����}��7�F,|>�Ӳ�	o*#Sp�k 8�1>��"M��<h�Vm�E�sӓ1̨��s={�9�+�𳷵�F#ґ6ƈqy0�4ZZ����H;��
6��-�Qɣ*q��wr��H`����\а��mw4:5��K�Ӓj�����c��H��XT�>�9�\��d$7'�ge<nLjG��YfI���`}}���ugFuQ�VX�&�/��ƺ�ϋwh� mh�`b��q<�&8� ����>\����F��`>8�/i����j�����@' 7+�+��ܼ2�R����/V5�=�s�QQH�K�X��\�d�[�k@a��y�';A�������,�9��F� }��M�����j?sh�lՇYu)A�'�+�,�À6M}α�#N�)]�w�����*����]��n�e#�9z3��Gjк�M�
��{��g��9%�1��{��%�L��J ����Z�Ӛ���\'kZ�=h~�o���V;>3�Z�Z�G'�1~��O�Q�M�,f�#���=�r�/�e� �S� 檉w��� ;��Cʫ|d*�b�,��y������]'\���J��"҃;Z��a�D�4��l^�{z$k��Ѭ\��%��*MQ�5G�_������%����s(���MIā�P��>u���[�6n���U������{�3���wn÷����^}�|�9�&�&��sC�-�p���A� N�᝹�E����W~��d�J\��T�`We��D�2�dB%BhK�>5��U#mm��h���HK�1h�i�#҈�~�q0�I��m��^n3����75�G��7he94q2˖Z �`�-���3�ھ/�j5#<�@8B��9���g5e��^j��\&����L�b@�&�c���Z�s͝`��Y�Ї ��|�w_�� �VC�֭[#m�����Y;�t��`�`�J_S��X�X`����1����������Wy����޼��_ի�k�U��4�Y�&@ ����1���	�8b&4cO8�?<1c��a�����$@��ZR����ګޫ���/9�_~���ze�����*Z�n��_�����/��;���9~�E�4�O,���K�گ"��r� Cƾ��ll�s��gr_���dhȼ���P+��W^�Dx�8>i~d���M)������f��j^[
#�I@�?m�R�z��@_��3x�@{��NpIg<ch1�.s���<�L@ʶI��@N��/�Ѿ,��n̫�!�"����L�B��9�$&@��Q`��������:���5����^�5`���-7K��\��A�^
6m�a�4GS�y��ơ��rp�8�$̻�1F�h�'�,��E�j(���L����&�~lϏ2���uZJ���}�4BZ�9��[#lm�q{m�5�jaw��!ˠ�i�3tσy�6�;u��9>�_�h{�;���������G�7?|�+W_���E���f��uM�Q���ͮJ�:����"�XKJ����&A=
	H4�����Li��zc�8�(�@T�QjրZ}V�JF�+9$� �� �����Ѝz}�]T�jL�0J�ƈy
F��eU4΃�sj�)�ә*
���R���x�G�I�Jը9���u/��1��3��]��-ջ��x�)e(�ٜe�M�޼������vZ�KR&��LJ�>]/�M+%����&���7������D�V5���,����$p�)��]�@G�$q���hw{�wh�	Y��l��2W��%&��4�G��<��k��x��!%�$si���s�b����	���QO��0-T�g��m)�O G �������eU9���\�-U�\���{�7�,��5w$*���W^�� *p��T]�W�XdL�8H���i�^9S��k��5��2!	�|��M|_�����6��3���P��4cd��^���˶��-�/����������R�k�/�� �S谳D�bZ� PR���u�8����}���oQ���W67���x�r��i�L�f���Ll÷:4Hss跺�XY���|��|�;17�@�����c{��[�[�_:���6vv���UDxq,j��g �G�.����,�?��?/����/������z���srn�̹I��,���TҀ�pP=�/�������O�a%�&�Mύ���	�J�b�5�01Fq�.��hǵ
*�:J3U�f��ec\N��r���\�}zs�1���;�ps��ƻ��M��bDV�/���j�"cJ�Lbx?Fg400S#"e9�@�k�n�fC����̀�=���f ?�T�LIK��"���`N@&��0��{�5�'�\aR�ĔJ�2�i���r)�-%q����Sx晧�X|�԰ٱh�og�W��4M���sî�.�DΈ|�����#?���xB��H���<(�~�+U�:#=��0�w~n�^�6Ȑp���R��\����͚L��4�QNp��K��x�f�̲ƨ=H�!��vFs�͇����ڙh��p�m�O��F��z����<RC�'/D$0�}������+۹h�
>C��k�o�Y��ͳa�}��L�=�	�G���>������a�a�"?ݩ9,O'L[j���!���ꕹS��0%0�z���2t�l�΢QKCQ�q������WL�v�������f5A-��{���p��|n3��,8�u;����a{���V��5��&��31�V��������iE�h�������3o������޾�u�pLbD�L���<��.���à�W�ڽ��T\Q(�ëC&0G�Sev�v�M�F�X�7�gJ�0I�n4D;`P���*��,�<_Gm~Y��n4� ����dck�h�,�2B�CfN��vG�m�sg������6R:����䝔,S��@^��۝qY�؄��������$(ɛ����_`*�&0�c�����E	G�PJÔDT�*^�C	�ו���˒f�z�r�PB$X	��>���]RYߤ�'����֙p���^������ň{D��8�n�A�NFa�(�Q��"d�c�u��{4ߞ�k.�#���XhO^jT����B@c�hK�U�y��+sFO�C$ՉY��c����E e���H�i�yR�M1!:����> w��5y�k�%r��ݴkh��%ߥ���=��;< �{]����h���������S%f�畫�MC$�e�_���OiJ�+�S�La�(�<�Z�da��Ba��|�Y.PsZ��3�ǃ9%tc��4�Լ���w�B��d��N����ה�)���:�j��Q�3]i2FZ��]��<��1���77����)�߾����2v[��������A(g=
�� ���XX�y������m��p܆������ޓ���O��7�[�GH�6ɤ�0E E8��s�r�K]E*+O(��1�f|pv?{��ʌ�c$c�ڃʝ`>t6"��mÔc�#��%��3�-�a�)=�%t��F}���~p�z������N�~m���2J��T���]#�`��a��b���pmٝ=�:�LTF����0,4.F9�QQ�1�0aʄ)�#��\ �C/��ל�$��i�s��*ν�{�$F�G������g����5� ��$A\���C{����S��:�) Wm���0�l׼��2�q	�a�!��T�V�9���&�O�ϼ��t�^���V�^��>��!T�_d�8�K`��R�ڹ�8��˔b�*�r&��h�Y��ӄ>�G�c�' �c�~1���0�O��q���o�i����=� �G�	��t�Q�~�w�U6jͳ��=��X��Ƭ��i��E%�{�·�Q���Ń9ۥ9�pdZ�D���7�a��M�IӉ6H�hư��Z�?U�|��f�!���t�[�6��'�7��q.���=Ϸ�}��+S敾'{�Pz5-sd�R�p� ���g�Ʃ�j�������o�`�x�"�yFM��{}ܼq��%�6�v-��ܡ,`>���)>I�t�e^�O�}��{������{8�������������^G%�6	����`>垃��w�ҡxՠ^��B�g �U[ZMKʰ��&��M?۠�dC��1��@#Aui�����c�^�v����V���h�4�1W�b&�`�>���;����.�*e���?��^*c$t^Yo�w���n��(B<
���G)�'��8�PE��iE3;����H�����7����R�!�W���' �s�"�^-;�X��`��k	TDk��Ā��$q�M^}eɰ�aq,�d��(t
2I���8
Ik���kO���3b>8o�E���Y
<�5BƔ�s�����(��	����NN����x�`x�H�9Gr���EZ��2�B�/���
Y����T�^������t�:_�||56���͕K��z��46�.f��}�@�Ș���K
�=C���y텘 /�K������ޘ�.r[��R�V�47�"����qr�o|�'LI`J�	�c���DS���q�L��A��yn    IDATL����XO�7A�M�[1���5Wd(X7��G^m�`|�)v����k�ylԪf6 �S꠆m@��&��tQ�̠YoXƷR��;��*��w��^KC��*��^o���.nܼ���"��2�6����	���cS���@<��ǣ>������y�ƚ�d��/~�3��������ӛ����Ɍ3g��ٵ�lZ�H(����~c���%�dd��M�MAΏae(�SJ^�.�i��L�;l�2V�á�����4�8��v�Љ���w-�-�q(mb�����X��bgo7�n����w�/G��K7-�G/wf`����!�� �����m��Ҭd�lL���G���&,��tP%]�.�+`���ʼt��P�P�i���"zgQRA�Ǳ \D�����9�t��X'�g�(B���W����o��&Ű.�I�A}Mf�	3���
\���Ҳ1>l��hi"�%V�n�!C�%���:k�j�� y�c�� H�IMb h��Ƹ�G�Dk��٠�o����ۡ����MS����${��G��^H��w��"�rS�1�l���%����.���������Wk��պ�y�9s+0�^ӻ�o�Q/�zA�k4z/����}^���5��z��eAΑ����,<���1��5e��!��K{�W�qj�1�;����lO��!�>b�V3�>�V�$��3��a��u�{��1Ӭcw�u���U�g�uY�F�:ga��$��u�?����o��$f,��vg�{@̬�u���A�;2� �'}`�L[����:T�d�:O�����С�c���\�~I�<˲�C�ԏ~�>����F���E)�W(%��1R����&@軗|�2��Q�v����������G�p�[��[]p��c�d�R��=���VP���֨`e����q���^;��3��j���bR�*��jMT�5��up���g��$F�
:Ч��}�+*{}����`p}�q	ʹ�A�o�����24�G�������nL�	=�c�U�~�=q�uI��-��� 9@ƿ��*	��>��D*$�jt�$?9��q��f���I�Q��H�U��[��R�&V)��3o���7��&�˶y�/C��O���h�U��U�j��z���Bb��UR�����k�����%�cF1�?e��=A�JJtD�q-8�s1O\:(�]�r=��s]�DSs�k\/I��[#sV�?wp=Sa^�t��;�/��b�B��bV�u^<�K�.P�`.�.�#1:G�+M#�s����t�A g�k�;�٘s�7�����C�"J�N��Os�~Rמ�~�}i�a���#ĴM�_n��1�ls3���255=�+]$�1f���[�Z�!�P�<x�����tk2��<��`���k��Y��1�;;�ti+O��Z!���?J�3T.1�k�����G�?�rp?Η
�ӟ��O�ϟ�����n;�PJ-��br��F���v�"��C�{'��\��=��0��ηo\&m;yn�.S����1C)=�y�Ϝ\��Ϣ:W��A�%W�=�dC��Z�x�J���.��s�wX)7�A��n߼�_�Z������<�~���8J1��i�QU:�mvQ��b�k��zX��a�!m���k�~p8Ƣd�%j\�L�ǪT�^��ڿ!��*�t�����׉�0�|��R��0)9��Ԇ$&>���^p�B)O(M}�@Nc
�,�����9�>�`�4�8\�`�=� ���Ԗ=.0,�7a��gv������=c�SNF֟܉�ש�%�s^8���I_(�sn���	��S2��W�����_S]3 ̽�%��=ك�� �`*i��)���4�~��s#&˫�u��}�8'�������{fA���b85�����"���3��\3���p^X�����P���~����L"����d �W�9�e&�JᑇC��T�r�kZ��:���|�����5�lOZbZ�A'8�rﵻ����&���-�����+����v;�"a�N#���������Z�!�����.Z�PcC�@Fa�<˺�Ο|��#�_�+0�G3����|�c�g�gO��ng�$�[�.�y1�k8�A�q(vM��'2:��#��D���oV�T�0�7%��!5����i�QZ���#8r���8΂��x���.�G=��U���Ȱ��3P��t�;�X��N=�kO;[�x�u���}�s���ByyΜ:�J�B�(q�{��z��E��C|k[�_�lVAi��uV����K�j�8xպ�.2:"�s��=cT�Wͩ�:���)���~�E��/�U���T�ROJJ�d<-A�`��*�#�H��؞r�O$�<��<�����/3U��+ A�`D)f��`.��﨧Aʠ籕�T&D�������}bGΝ��sS��|z�`�:����	PLJW�ϲ扪4\W&��KB�v���R ׁ����=�'%x�#���$57�^�C3C�w��D1�|�?a�(�T���KZ��K�k/Uk^tM������cU���YҾ-2ꟀUL�g.ن�s19s2�D9��Ʉ��9��L��g��$�����y�>���g���y�O0����5��3c��2�#��y�"�#m���"���^+8����x�p�p�om`w��4� Ye����'��VW!8[M�Z}�^��������S0�0��y57�Z�I8��q�q��:s�菜�o�#�ʾ��}I$�7v�?�+��>���~���\kN��Fw� ��D?���y@�*ኧ�DUڈ\^[���2$E&���2�^BeyG�?�ƑE�k���3B4 ���0������<�wb9�y8�^���G��U�?�tL����q���,�s5��%K"S���xh���(W"��Pm���Mp���#�좙ѻ=؋����1�Bn��")]H�Vs�,/i��/y$=S [����d^"R<���C�_SO�x�O�>m�)�&&�ϓ ��1���aN[��Vv�	�OB���U����#����j�Tx�?��e��_E_sɈL�$s��ԯlS�'&��[�N
$x���"�3/}N�(5���V�yf��x�T�s>���	�L���_�t��8���� I��+f��)U�iԊ��@L���?Y�w��2M�̝a?�E@��� &M8�3�פx��^�3�Pt�ާ�-��Α$k��{���[�w��;g�W�����,Y8�?�[	�����dvC�;���(g�<��7sY	�]
f�M`��Yqyl6g���cѥ��Y
}��QBDg]0���sM��
���7��7ol`mu�;�#&�*㻿����ןK��Y��{�1V�6q�ֺ�9CնvZ�GV|�>2�De��0�vO9���߿�ﾮQ�u�%s�e��/짞z�����6��l֭��������R�Wsy��ġ�����t ������9㷍�2T(cXO��*OE���j�6�L���?DƂ���T�wwv0�Pb�p���X�������5Sg�/­�\�}����lۭ=̥5������n��3T{c��Fh�x����Q��:�X� W3˦�AX�>O�4_I&����;�� �m�oQ{�I�Z�Ck@�¿	"�+	s�{ə��	0�P�W� ��9�NJ��ҟ$Ŋ�ˣ; A��T��lݙ��r�O�o	��Ȅ�L*<�1*b������u͕�Hx���\��OLM!���W������3��;�������y����c��׀�w����R�%U�H�en(��L���KJ�jvO�4W���k�^DՎޣ�/�X���L���KZ3N�x��W'f�\��w�ӛ�Vm�	�f���-[�/�+Ǿ�`��/�+��攨u�L���g�Ü�|%ec�L��j9LiGnN����c󞃹��S��@�}��W�6��VA�0��q�=w�om��'�j�s����ߎW>ri�Y����ls����굛X>t{�6���'`�so�{V臅�H={�����塇V�EE�$�# �zh�%�K�6O�܇����[:�!s�F�(���i�9⠪�RI�(�@�X%x#��)��F�����#��Q����2��Ge!�j,��b�\Ř%;=�u;��*�������6�Q	+�9<r�Y��x��'����.��1�����25k��8)�ӎ�P�P���lai��.�1ֿ���u���'��^�*m�Ȃwf����f(����H4��#���^<�{�i��Lis�{��O��q��Y��"8�9��%���KP�D)�9�F��}l�c�q���ΒSg(�ë<dD�0O�=�X֛&� �5��u��Hl�NBI��-����s������<�&#�>�H߃�c�x�͋�E��,�yU����	�n�jgp��*\�BI���\����@� ���aq���5/M�L�	4u����Z^���k���x�A4I@ 204���uC�=���pb2S���f���g���H����;�~d�C$H+d9TS��ٴs��za|�1l�n(&}?� ��Yl�s�K��b(�' a�!o1�q(<T�����Ii�Ơ��g/b�Y���|����7��o{�z�:k`0�M����m\�z�������A��G)	� �%h}�p0绖����+O��cQ����%�.�^�У��_���n?��܂e�W-�VD0��+8��� �_o�A�R�?�>4��#0Y�p�2%�l�~<D��a�TC��V�?c���lu:��Ҫ5�����6�BJ���q�3�x��)�ʗ�6���o_Avx7�{��	%��0.c���1���,	L\KQE�Y	�Y�˟y�����A�~/�al<�2��ڸr[��|-�w(� 0��Q6t^�4����&0��S��[��Y�1W\�%ȸqc�Ժ����I��$N*�*i��D�"Zњ`���_���Ke�'���@�%yڄI,	�\c��R-���W�K>��.�к�\����aH��΃=����x&u*��a4�˽�Y2���ǿy]ah�շ�>��D�~hyш;� 0b?��m�2�x;�A6s?�S�Q��k�-��.@�X5W�G�l���_����z��,��)��Щ��$�,�wȶ�k:'�鑙�}�̰����ҋW�
�|�A\�p����IJ�|���}�3#�&�sr�j�Pb�ScC�����f��n�lo�y�������l��1 |��������E���:�Iw:!�cqqk�0��4Feg�c�eGEkw����߆7��<k��Q��cˌI�����W�cvn̀���6�v�Ay�F%��F5�&},.4~�����_\��_F8nC}I��Ͽx���O|����W0���dm��j�e.b촜fQ��&Q��&0�Tz�y�Th^�7.��$��qS[�7`7#Z���٣����s��K��eT�{�6ۻf_���2��jKY�>})b<��p����[��Ǯ=�����!z�!��)N���^�W����յU���2U<K�V%4nwq���P��(g�����ܡ�4/5�{�����׫y��"rb�>�}m�t��ã��c&+�IH�V�4�I�$<����7B�C�$II��.�+���^g�c?�Mk��׈�p`�D�S�s?�Y*q�S��<�����*m�4�;���䜲�Pe�#�~
$�5P�$+ �&ͽ��f�	ɩ�N����Y�vF~�K��QjZ)Я��F=X{���s&�L��Rk���ۇ�����:͕��ϧG^�׸�c۔Q�΀�/fl2�.ъg��r�V���i8�c���0�C���2bt��	�Z,U��~Q�#�isg��MX|��A&kP�r��Y��֭U�{�=���%��Pp�.@�l��f0eK�Ͱ��%2ڌ��2�<�Q����*��)O�E&�\-�v`y��%k:y�>3�]z�"��Mo�_��W�����G��	��x���P�ΡZ������m��_I�u����+Q��x�z5��W���4����{0����7��G>����WW�xĩT.�yH�:���V��\��uXD�DƵ�����J��8�A2B/��iF(�wK�Y���zKi��l9�Y#mo���^�	�=<p�4����ۛXk����ן�37� +�T�L,s����O=������M���t0�y��x��u M�(U1ۍ�\����ϣ<��#��%P`�<}�t��\�'�"J�W*y=祴����\�cK�AK��/P�{ȩS����ad� F�8g�'�xU7�mR�8���'��������מ����Q�\�*��K���Ȅ�D@G1B������#�#������$1Y͹�ڋ̈�K�zu&�K���41/�y�C0y]1���&��s�͟)޺��j�?_uv�s-���L���5_���k>9���F{� '1{b&4�WQ��w���Z����gXＤh�ڃ�o�Φ1���-�{��l���X��4SR�y��&�;���JD�7�%M��w��]��x銝�������GOX[�����s;[��Z�4Ph�m�M0�b�j6�t�:;�N��H�~�e�r�Q�֌��|�*�p���7!��X^�����dX�<\~�
"��5f����.�����P��WbG#)�V�Ͻ��S�.�(��n�%���3O|ӯ��~��F��h��S�q� ��	D%$���s�a�[����^�*0����T�A�舒Y�,;Q�Z��R���̝Y1	�`~�ڰ���)�i[�as�	U�:=�\<��?@��1Ǡ�~�r	Y7:��FO��0�
�x��}8�xO�	{�GN�D��SO~��ñ�J�;��z��|	�^��(F��C!��x�����xB�{<h���DR�+�H�㘿�KP�2�ʘ��p���t�e�#�%����^T�ss�aҙ�{W�N�m�=��M�K���VDy��'�ỨfW5i䨧Ը$r$��O�,nb4fI�^��<�~���փ�	��ZI��\��V'��m���E���)����&����ك�dO���;�܄��������׸���̆gH�_��4E��3O�<c���J!��Np��ߙw��9�g�#�{Ƙ3?;�ʽAIV	��]e}y�۳����
�$!&�g������6����������E��톊yt'���ek��.U������,"��C(�ج�QN��#8�����O �2V���膲��V��?�>��?s�����/2��	&�<yNw�8'}4f汶���`�U`N!��p^U�Z�����WV�/}]#�=��K����}�o����ۭ���q�L��\k�J�M�7/2!V.���<�L���A�&y�8�/$j6,��R)�ݨ�Ѯ'�ב�:�ڑyS�7kU�5�P���\��1z�geC�W�T�����Vo���$i�Z	[�;��J�Yoki��W��5��G���s�n��~��i4�,��{�ݖe~�f�Cl<si&���j`8_y��'��O��V�~8.�ً�	������}^ ���kMh3Q��O�l2�MNS^WwH�8"�	H0?O+���A�R͉�H{�j���k2R��h��XL���U�"n���E�V��D1�#�.W�g�Z�(�>��sb*�������ݤh?���׫�=�9�Cy>	��ob潟���2��A�,���{f�s-<}P;zq����z�¿+�=��gh<S���1��*�}Of��_�SO=e��DNP�~�l�B"�v{ϴB|�Ѩ�TLm����my���͗⩧��c�=f5��/�6�-:��X���9Օ�kմ��QH?+M'��a���7	K��Y�C�#:�2*)���J��'�x�?�%�9}����@�f�5�Uw��
)Z{m��mbfnw�v�Y�D]i�C��^��J9�|���<~��G� /���|I��#����o����,f�M�i�9�H2/��4���L�Aܹվu���c�V+�J���c�%�H8��l�j�Q����sq��r�RP���v��,�xÃ�������=i	h�r7�;��d���+�=>G    IDAT,�G)�Dco;z��󸱵�?��cA+��z�kP^��G�P�k�V�a�����!v_���01;zm\F��1�9�(�@T�K͋ Sk���9"XEP�{"�{x�K%�[ ��E£�
T�W�g�#լ �`~���="��'�^���&���V��R�ݞi����Wnv�|�nU��4	�zH.fJ��1y�[s�~L �"��V�[�(���\>��7�\̘?_ؙ���+�����z�b �$�5.�4x�j}wO<�������o�ݨ����Ik �M�Ud|Ú'^�H��`yO�k��}���s�)�'�|�ڠ����z�s��-�k�v'Y�6�k�������7o޶�vw[��W]�Y��0�����`��6C�&J�by��)��V�Cop�+� E!�u�/3cr|�ۻ��y"�'Y?�w ��5fYE�Z�s�����q��-�/���m�z��1�y��R4^=u���Μl���5�ރ��s0ϲ,�������|�:�&���j��Z����RtX�c���=��8�DJ��[t�>)Ғ��$����Z	8>��C̕M���ތ4�2*U4��jנ�A�7�+N�Ee��_x���ADLC:����w�=Kq�׬Tp�Rǹ��Vg.�G����;��[\@R)�k/�zw���Y��Ec���V1�UP鎑c�?b�����R��*0�Ҳ$YZIi~~���!�Fĭ��T��\�Dߧ�}�����3U�B&d��Z[I�lO6�	�f�cI�r�]ҝ�"�(���$iiT}M����t��gE�a�:T��ZҔ$a��5���K�ɉ�l��!4M��?�@y]̒�:'~�=�09G������_Z�7Y���\<��!8hNՎ�,���h��7iE�ԩo����՞ք׹��GE�D���j:֠NW[�G&�m�|/Zƽ�{Ξ=;�%�!�J"���{o�T�#A���*RVBf>���eW�B_�x��1�(m^�$N�,0��������*�]�it3�=�L��0W�G�gŞe��;}J�w�����߾�jf�oF8�4�FF�|�:�W�����N߮�������7<���`�s���w���/����n���,���~��?��g�I���f�����!���F�������:�����î90���C�C	Qڌ��1���c�(�^�x!�vַ\��q���^I��#���t�_=��|��߼�o|�[���eXV����c��o�9��-WY�;�Lg�z8v�(��M�>d�S���3��uÙ�|I�U�N�;]�=qh��c�(���S����Hi~2"R<�H
�E �(x���0
�Q�`�w�~I@�%��U#6$>K��z�LZI��AuA��w9�{	�K�����=l������ �O���*��ݟ�V������S*͏�+��"�M��4O�1%����3�����Ms��U���ϣ�
1DE)ݟG��=��[1Rb(��,2��.�>H л�����-i(���
�RL~��#^��J��W{Y���� �������p+���`)_�K�v躝i|d�"�["�jP�sn�i�\�k��H�� �cTH����k��g¤��E�S~c��"HL}m�i� ��^oNR$��dXY��A(2M �V�!smm��cv�������͠����J�jO�G.]����G�w�=��R�Ê+��Q/����ǎ-��_�Y��9�3/��������_�G�cBN�y,������ͥ;�)��ѧHT�d���+7������N`��Q��U`*�ґT�E�T�樋~42/�
�	�I����2<x�>̤)�+u�mn�6��'���O?�Va�R4+lw�Rk`9I�H*���@{�G;6�mtYδ�b#ĥ
����;عxQ��UX��U���#�&I\DU�J\� ��@��%�=.�b���eN��K�b�HXH�dX���]S5q�^����|��H���9�6��E`�S�W�.�l6��ÿ%mH��=bHD��4�v.i�Mɖȿ�_���r�S��G� X��g������f��\��wj��I�5��Ť(Ӟs^ꓴ*~�h�z�k�ؾ�hh؎T��+@�̣��K��=�{��W�=���O��� W|��甧���=>]��x�>�ϔԚh}��D��N����l�Y��dƾR�e�eZҹ��u���V.5�|U*�vo�Q�������+d���Ŕ�X�`�#��]�
$�Pޕ �kS)�:�b(��3;i�nL��ghW�|R�������w����J���%D,rhZ�/�p��|sc{��������x``n��n�E����#�x���EQ��2��s0���������녋���j����cF��E(���x�<�/b"/w����u�m�;e�@�M7"�s��h�A� =:���
�C\�l�>�z���}��E��Ra�\C��%8w�9��}s��B��%����s;�T�����ǹtoz�P	F�`�����:>�����+���-'�$Ҥ������7P���t��*�tP͂i�&V�E #�����湨B�ږ�^��4p�4���`�>x�C�6�`cj��jL����'�Zs�SjO�/�'�O@d��������HNM:�W�$i���gJ�@/�+��$.�^붏��W #�ϵg�����0W��7/	z������Y���`?=�����;����|��������,������R�����1�<�����sQ<E��q���}/>o�7~�I����cIc�M9�.���L���Ci��軩��#T�;�����d�1c{*���v�,0̌%��	?F�6s>G&�����~�a�5��
�s�T��\o"T�/�_~E]۟�_pxeż��:�ỿ����ox5��Q<20/WJ���4�x��QoΣ�ccs��3I��!�w��H�j�z4��b�'^��c?E����m���Yd����G���|'��TIma�
qt?�{�%�0�"�b��{�f1��b���gMkrz�Ȋ����v�*G��M�H&C���L���p�Í9�G@g}��C���ܼ�v�����X>��'�]�Z��A�f��$5���+gPp���I��+V��	e��E�f��C�U��n�z���]�6�̳���x� ��dҨ��D��EH=�@z@�{гZ
�U��v��{q������?8��h�Zoݧ��s~�
RD��uDM#�W���%��3��=�yp�؋*Xͣ"|��k2H;��\ ��t�~O�\3��ԃ�4+��ճ�xͯ��P_�������$e�WZ	�?�W��Y� ���`���1Z�gjx�{i��7�I׵w=�r�q�$�|.�i�-��c,�Ȳ��	�\�/�vm�_ -���ۓ
jFʩ1�����켽K���������C)%&5ӑΘ�8d���XN����=�,�������ۛ���s�v&�QZ`�{�cE�^��?�㯿�x��߄2k$$�}`�l4q�⋨�f1����6B�1A�j�Y`c����7����ff�տ���3p�����/��+���E(��	�33ɝ��*$������w�"��;��f�9~���!�z��ꗏ��H�-�y�v����� �L���a&+�Xc���ju\�}���q��1t�\Y��a��>1X��D�5��S����x��3X^\D�;���'P;}��D��~�a�rz���obv;C��.j�1��>���=�"")�,�փ$����N�!�\�XzۼR+�50�V�������%sփ@��߃���4�	pE�/���8�<���)�лD4�{�}��J��+&��Lf�#�/��	)��e�?hk�C����w�-u����"�T��� �{�5�vQ#��bv4n~�$Y�=$F��k���
���"�����{0/�C��c�g�K�E�8�� /	܋g��M��*q��`N�6��q��4�lK@N	X�������G4���H�ّ㥃���Ա�5ݰ��f�=3�@7�����6IS�����;�}�Li]�|��H��!r�6����;��r�8[�2��z�.꤭���\�!J*V��xl������m&Q0�1�L�Y�Ӈ8����B��}S�\2��;���?z���;z�x�T�{0��TH��蔀O��\�Y���_�rnpƍ�!�f��ڗ0�F� �
�J8�6P������;��g�r��Wq�Yƶ��w�����ѫ�0q�d�!V3x������M��S_4g�E���+�^�������j�*,�#��� ׷�\��|T��z�)��NO� �zB��Z6͛��<��QT[Z/a��J��{H@up��_�,�}_<���V\q�=�x".P��L����K�T�{�.�Ps�%����p�4�E�rT��vY1 b�D���ծ��e�����q)2yI�Ź�z���3���S@�5��P�7%������t�E����I�rFԺz&�H/�̾ޭ��Z
��5o~}���.���(�Q��%s�9�C=u�.��Z�@ɿ��
���$󲩷�P�W�J���MƦ��9s挩��1��v��c�f:Q�����鳈}B^���bW��(I&��L���]1�*W�6�dT:�-�������D��ʥ5]P)� �M���2������"c�hXw9I<�Wk���;���#����e�������y�џ��n��}�`�R��M��
b%����_5��$���T7}�x��<w�AR��F�:H��,�ү��y,�;��}G��ݱ{�Y��,�R\��ǐ���_©󧱸��g.]ĉ���������MK��$�Y���j�Whe���7QK��܃h�f��~7v7���< 3��y�*�C����50{yZm`�ݲ҄�\G� ��@�� zp�d��/����rB��`.��� �j�$�%\T�ÌR@���K��b(<Q<H��`aD.	��p�A�p��rS�g.ش^���-p�5����W�\d��^f���F����$�N.5i�=c����y� ���^b�8����O�eQb-2���g�?Z����
��ӻ��׺{��Hc�'�=~�$�����p�K�.�v��x��T��#9J�F�s �<r�;��jw^g2?��4ѷ�d(PXe�noc^t�9��y�(����v�ΚiJ��0M+���������"s�~�َ���7v�O�o~Ƿ ��H+tN�"cF�,25��v�R�R2�tz&�3��~TZ�!���ʣ��}���/��1�̿p��O���>���~�h\B%m`v��R��Tf�P����ZQB���� ���;6e�+J8"F�!�>��=J2��z���j'1w�P/���QK�H�:8�6q�����ڽ.�3x�K_�(�p��Y|��ǰ�0'�Ød�!J��k��d�%%[Xı�eܸu7VQ_�Gw���K+�m��q�W�Q�b~��僢J{��I��#��e��J�6c�"�y�/���\�_8B>���<�REz��Dh���
���:���j���$�A�}��ɿ��v|�'�Z{�=ҝ �-��9��U����_�Eb��9ȳ�T#7���%��DRҤ��<�j]5Gy�}[���RJ����ȟ#1J��[z^������.E)X�k�x_����T�}�N�y���CX�4�ի�����Vh����9��ז�ooJ��ǃaf6q��R�Rz��ۥ�]������Xb����n�U���̩�=$�`�79u��Lm��2
��E�O0���j�W�y�Z�eK	���N0�׹7AHSG��v�F����'�����b3��͚L�qܾ�nY��V����h'S��!�s|IDG���Oy���s�8�>�e�v�������W>�яx}��H�
���}`Nɼ(y����'�E���+n�I�O\�?L0�0��4�I��~y��l��*fΟ@zxΤs��jM��#�X:d�7.]����ϟ��=���'���%ÒT-�+�L}Ī@�6j#X"�d̪EC�ӲyVϔ�A_���a>��u�6��a`��-6��+�Y2�a��
dL���1͍���ɼ��^���0� Y�w��*LJ�p�W����j݋�["(���Ҩt3!	؈�8��{��Ty�l/E���qJ��"Rb�]�q�1���*	��<��yB�S��1yfï�1s��t�^b,����\������e���Ns~7��>���^��ڋ��αƭ���z���^`��}L^>@�$X�S�}b��C����T���J C镕�8��ο��`���ݮ�����^ꜻ��=�Gm��'�O��B;KKf�g��`��1S��4op`����L��3q:��͊�􍉘�]���~˫�Z��܌�E+�Ҩ�©���Q���R>�H�n�礆��nc��sƭ�/�{!t ��<K���ݳ�W��ٳ���e��u������o����ڣ���Q\E���\�̆��T�<�!	��lb��x�"w�C%Id!q�i�`ic�0V�9�y(�8� �*��J'�8y�b��.j��3Q��=T�)�ۚsU<����wVQ^��^�k^��Q�*mQ���W0�t0�TQ�KV�u�u;V/�>L�ws�h__G��1*!n�Di�<㓼l��;?,d$Y�{1��=�i�����+K#��i�QIj�O���㉧I��=�� [
�"�`�;��ᜳ�$b:$z"�_�v0�9���Usi*̼�����gf�.���;�QҒz�K�^������N4#��5�^���p��.�?W~�=��Aѻ�N�nI��|��.�� ��=�����s?/Z'i��{L� >#��i΋�}s���3I�
�Bo�x�t?F�n`~g�;��	獦�׼�5���+N����s����I粠�d�Րj���B9Ri'�;��`Ksz�K2���9�CY�����1����,�q5���ju+���϶NL���~>�w�o�:lmo`n��#�5����*��Ǩ�#��I�i�;�]��#�N��|{{tZ�(����%�{�@6�N�>�c��.������瞃�o��c��������p"˹��Y��V�(�!)��l�*�!@�ң��t@���,�&p��fږ�&:Qݑ�$A�
�RN�D�Gc��@o����y̞ZA'a0`�똽,��:�$�1����v�]h��U1��34�)R:�0��*����	���u�����εUtWw��G��R�4S�`���v^S�)���P&b-¡9�*n#��Ph���`/0(-���f������9k-H�H��"Ȍ՞н�X��j�x���|1)��#I��"��3ϼ�>yi�	��>�3�7I����y�X���v�B.�Tt����Q����%��$L���N1	1���9��|E͈Θ����ʯ�D ]d��{^��?S�����Wkƚ
~�0�W�X�����8p�	�'�"��~�H+��^�1���.���(Ef�󷽽�7nb�ʙ�xm���^�:KZC�&��XM�Vˤ^�#��`;|N�k���K��F@V�|�A/����t�ƨR[�X�T�s�OG����v����d�XЩ/Llb�>H'� �1��p��R������pxy�l椏�&��w�pgciu��뻖��Q<�a��P��r��K<����|�+�} ��P��e��`����s���_�����e�L��
��yRqޒr�9����TZAID�xD\	�!�QHW(�,�#0�m7P�bx!�x 1���0���?|��,6��{��8:�Iܨ6&ﵘ�0"�Ҫ�I��5'%�,H��aL�9�ȔK�[�
ƻ=l�x[�oc��A��i%���HD��#���%��Z�W㉈i�a��T�E�Ef�H|=��L��4㚽�z���Қ��E�2"�b� ��m^��IpsI`�`��|�;�q�G�__I����h��{��w�ӼÔ��ja�P�:ݞ	���_���}ρ�1z��6_��������&��Ҳ�#�[s.���:#S`    IDAT��f4�l��ÛX<����} I��Z܏�����
>O���x��ă������Α�_&x�����ϟ�Mc��D47�������J��A;л*���7�i�R���|�`����Ŝ�r@f��]���M�`��jv1k*Ĥ1�C����Z!�hk ��$~���^��>?�h}�����?�s��f[��x��z����{ph���r��)�%�C��ma{w��"����<�n����C�$�_�XZ���3������� �����~裟��������~4�X�
s�ΰnb�T��0������W�f�VP@�n�7�MϿy�[e�8������0lg�aL�T��fk�6n��ox5��JK��)_+�;�}�����מR���`��bif�T�LK�Z�_��,~8�aH�<)���a���^����˻�KH��n������\�቙���#O�dFh�\���{��D<�6ic8�I��"�bD%�{�}#�53^�*�6�J��9e�t�/����ޗKl�N�H����/�G�%CO��|�}��.P�#�&1;��h�\4l�ʫr�9��u՞��@m�k���#iY�iu�h������,iy0d;w���*2TQ������ÚN�_�>h�m���@k�ݔ�z@�k�����@>T-��9�u��4������XI�l���G�I�A2�@�Ǿ��Oi�4�t��5�٩5�8�[�,h�8��o0ݨ���Ԭc���,���na~�@��j�E��^�'P��'N�@g��D�GVf�e�ԚF/Yǂv���;huڨU�1Ǹ��m~Gs��YZeD�Mc���g�<��}�[iF���^#�׾�{
�Y�U~�ß�>����@��J�rxi�Z=E�.��l#^��Ln�^���ͦ��2P��ˍK '�������M�7�T�v�r۬?􁛛�8�9�F`�k��̻����w���?r1����h�f���(A������a�ް04�z��a^���@��p�E����v�}{��װy{qg��(A�#�%:x�� p� � 9@ƿt�c��$T$�hN���X �q�=!;�	�fӾ�>������`+ ���_�V�P=؋�ӻ��T�űr_Hj�R�$J#0���hn�D��@�6QO�=h�|��|�b���c_4wR��6 "b�����/�\���̞��AX�7��? 1��!�W뤶��,�u& ��ћd�3[�s���ѓM����ń�Z}d�������	�p��@�?�_�&���?�4�A�@M0'm�7;�:�Q�%]�sl�{V@e��?h^g�8Ə���F)H�����h��پ��ǹ� 	����u�'[�<)N���Q2G/�������^j�8ƙW�J�.~�ߋ�������|s��VJ�v�jv�~I\����D?!)����[�K*13���gϞ>�ޕ��ů=̾4=��`~�V��ŏ����O�۝1�YH�_�"&��Nl��I8��!7���F����Xlnr9�����9� ��R2�;!�y��?��7	2�H�y��!ΗL��[�Qo6p��Q���quk�玡�<�Ƒ%$�u����1C�h�z��UT��`������0��G�IV����ظ���zY��F���8�p��h�Q�a��"�L�`�3�r�@("�%{�<�u�E��d,�d. *J^��.���E�������LM$��>�G�����!iU�j�݋ē�ez(hlFi����w/��TYK1��
�<��K
�v���<H%����n��x"�:������A����Iк��6�k���̔�Z�˃�9�]�O
�������W������7����a�&�gx�.�{��]�sQs�w��T����"#�����D���V���-�:=�(�ox�I��kʦ&)��A����]>�~�k>u��fWw��I�Q��ɹ���]��=�=ƚ�)	���g�s��h�7�S��`�8��	��͎^?���k^u?���1[o�R�g�[�vj �q	Y\��[�qBA��)
5ԸMm���mT�8u��?���K�_���S0g���~�W�������Pڌ�F��P�R9K�E!= �=�p�QM���	���f�''+�a����;y��Y}����t��0�ښ��lA��X�cak'�;��x���66�>⥆9��]B�Y���LȎ�&p�l�Q�|�	6�Lk�N>�����ڍ[������&�}�R�q�
�̕0���H�!!;��3�X�f�a4�:�H�&�T���Y�פ�nR�oK������jv��ge�"�ZSI.���3O���R����V���b���	��W3͓lު�.M �R�j������2I��+[}�Y�	>��u�%#�������m�|֫�siO��"@�u��[gX��Hz�e߆.l����w~������"#^\�"c����Z�D��g��;���xfĈh�=�{�>O��T�!��g�[�f'�heK眈0�}8� �[`[����y&�Ȑ���'6x��,�`p��_Lk}�^B��О�����{��]p�����֖{����O����w���߀������\S ��GX[�m4jĄc���b~�>�x`eP{G�#mݩi��z�����?sr��_{�}izpO�����̯�������!�	V�l�Q�UL�BtƙK��lU�Rr3K"�*J��7�Si���E{�ޔ*�'bo�`�L<U2���{g40�
f1��:���ٵ4���,ת��wp��gak�.�u��jh�4P��A�p	�?s�!�Nϒ��wZV�l��o�!,�[<�ё��X�M�jb��n���;�qDdȕJ������<Dh�(�p"J^
�w�S1�P��mIw��_�������f����_�	����(7%�:>i��m/�y�����0��z���7�FB��K3��O�� ��'3+{�I�Q�;1M~ν��wz����(�����@;e �&�"�O��e����R}{��ާ9� ����(���xf�3,��s���8��"�\�}���w� HVdR���b?�ѥܷ��HPk��K��ж��H����c��NH�F)����ٓ	�����]^9b��m[��n'�>%�K�����m�e�K2��	BӸRk:_ %e�I�F=E=�������=�5nܼj4�s���&�]��"J��>P��ǝ�]K-;�B���`%��9��֫�ͣ���g~�ү�[�)�_��>�?��?��󗿩?L��*h4j&����I�\I���/7���6t�;pCr��0�sQ��߹��7���9��:��;#8���c���צ�?�]L	y������V��ԙ�p��u\^��v4B��"N�;���-��	���"�f�H�UϘ���EyY�T�w9�,l��z#�����X�`C4B�C�,�����F~`��˫���y�k�/މ
�y����"����K!���Ǳ-E"�dx�q+��ߥ*'3&���s���)Zs��m��oN\���1i�$���~����Kܑ3XEU��ȹ����b䍉�����^/1��Kd�t><hhOx�\k������g�s�Ao�{�pR�Ե�ĸx@�{���>�roo͝W�QC�T�z��@/-���g2��xM̅��3�T�^��(���Ϗ�վ����YK��׾֊�P2�,l�P��{E{�?�"�U�i����2�]�G����>}�K˓PI���۶}�}j��<�+��#>efm/���08���F��s�k�E�6p�<��4Ei���^�0���y�n_3H�]��P�F�|�
J�t�h�.a��6:����i;Ff�ɓh1�&CT+�>v|�G�?w����0�������ӗ6O��O}�Cׯ��U`>3�0�7�ٙZ���� ID���67	���rS�<�}��p&&��8PnzJ�p�T#a�6�@W.!*�d��j%Ek{�V�ꟽNk��4�xh�h���4����CX��4f%�p�Y4elY���G���5�Rl�@������I�h˧s��%F`%��!.�$��s�E 9H�J�<O��L�����^��
��^�$�l��	WdJCR�
P��T�u�w}h~����}V/Qy@񖴨6����鉸T���{paIVI:�a���5�jV�q��3G^k���3S1mz�g����3l��И�J��3��
���������9|i<p�.��h��S~���;��b�\�^����"^��W�#@ˇH`��R2��LEX�n�%��9����M����Q�۵Lp���x�h)�9�-f�λi0}���s�^��B�Bh�g��9��K��^��^�p��<~���!v�7̇��τ��o\Ɛ�4���o���`�1�kb`�w�����?Q����������+�&��i
��W�&o��`����?���|����7�G��K,a���`N��qXy�/�^�L�����_�<m0L�/b�߸���d�*R��9�܈�(H�:,�+��M:,W�F2wp��T�	PiT���&	D��-_|��2��k��CsI��fls���=�MS@��<�#s��a	�@�	�L�AԈ�U
wxb}7) p��mΝͼH�$w�>����'�z^�]R��sب�'�}�6D\��
�����A�1�z�D����b�|l��A�8e�筀[�=؊��56I��<�O "�A�����,T�o˃�΃�g�����K�z��\l���LR�~�O�/�|�_E �[{���|xƤ�G>Wd��=�wO���J�(;�T�'O�&u�>���1�^�}Kɜ�!-d[2;�w��7	p,rBc�ǏǱc'r������p��i�f1G������L��<�"%v���,d���G)��� LE8<��5�Ѹ�q`f�f5h��^�����М]��V{�UX#���e�/�@�����i9���ܿ|�#G��(��ŵ��������O�|�'������jde�����	�y)B��]Vroz(�h�o�N�b��s�δe�-8c�[��O�5�N�.78C5��F� �t��aa{�J)E�ɭ�����TJ̤��BO��<�t���40�NNf�q���HM�$2-��|���s���o��1�����#�����}jEW� @ќ{��3%bS�>0C^�+������)H)[�7T�1�	�T��A:(2!�$��T��՗�3�9�����>���m$��v���=$Z�G�ģ�Dy���.�H�s�����������Ewu�������1�5:h��}����n�wqy�=5�.�oiO9�jF�Ȥ#m ����c�0�ؕ�}�K��%�}u�r�(N�<��u s��ё\sE�9��u�/�W�IM&]}�(�U�,W��2���-fB5�|q��c�M�%��3��{�|���^U�v�J`��,����`Ƹ�<=mGw�g����tτ��m�6��`��1B�$� J[I*�J������̉��e��W>����/�e����s�w�3*�XS~��?$�����]rbBri��g~�>S&;&��i)�R(�5�VE���O�%�`�Nvejz����s�G&'c�����ǞS0��������O�Y.^�g\ǧ&�0��40�"�X1��Z�4�x����	@we0b��F�~X�g~Q�dB�͐1��@�nϪ�!���d�L��d\���0������>��i4�f�{(�b&d5��Cy[���8p�Z	�f1���g��Νn�PL��E͸8��D�A`��D�A��̷0�5X ��xNo�V�D�t��<�.h��U���M�!n�z�O���s@+ J[.�ޟ�~k�HD3~$�r�B[���	2\�^T3���P#��Ώ^'���A����6��a��-s*n7o���c�9;{~օ������{�=�c¨k�7�&~��]��3���5�קb�"�a|�j�-�`�=�k����G��g�"��z�y����u���&s�A37A6�]��6�	���6�iv4��hf����P��Q�����kK�]��Wd��4*�2�Az��çOhfS~lZ��Zi���t��VE�`:�܄c����T����y�|>v��
Џg��̯����|��/���Z��x"+�lF�.���K��5f+}+����z���^(�&E&�j7��f	�v�lY�Y*፿
:ԫ�㎍�X*'k�+�(���`,�֞���{l�ə�Ga��z��nM]L(� �՟�y0�+sa�N��Q��%���L��%C�����3G|�Ψ�մ<#%��3�P4����.�P/�ךڵ&� 30+�� ��b!�`�h]�u��՞okU�(��u�����~x@�2�(�l3e([[�F�v`��"}{��=
6Þ��5�k������v��u��`�A�l��F��DA�V9��Ycbn�c�z�:F�[-K[h#���i�s<LX�3l���{Ĝ�`��H�߹�h?�s���P*T;�X�9 sh��aC��9�<09V�.����=ԏ�g�S>'��hчn�
���J���L��d����0��
ޙ��?�`����ݒ^�*׼�Mr��~������fv��յ%9y�LM/(���1YY[�����}͵���@U�M���Md���=o������>윂�7�y�U�~���^ޛL�$�I[!�4 	����� hv��@�~"���4��r|W(l(� a�b�0��R-���0���ċ�r5�R2�j��Μ��R��+Ҩ5�R,��];�[�5�/K2�ع�ҩFw�pf�Jݓx`"0g�8B�&���N0�m|�$ژ�z��B�����`3P�F��0�k_�q`�߼��;
򺙂��3A����d:m+ዹ�:�P�^�k`D<�@�k�*�1�w6��̣@���!2`�*��
p��	�}��cB�I˗5�R$�r������6��	+:���X ����G:*���> l��{��c�_��AQ �nͶ�ǁ���?�������{�"���m^��Z��w��a���y睧<�(���PT��#���Ϸ:�~O
r* t��s| ���Uk����u�B�sQ�bY,�����E�|xbbR�3K�2���1u���V:%�d[~����\q��Je���R0�/������ݒ�OH�7"˫+
�J��5�J-�=m��K�~p�η��d�x���O��s
�_�ڍW���|��6�;ә|_3O${
�`F��Mb���X#�	��v��d��q�G��8��dG�g +��H8�wl%@��b�<����{a �d6m��jə3g��˫��V��9�8w��i�s���h�(-K�b<�O����2��5��z!8΄��V��DJm�����L����@�&��&p�-db<g�&���7��<b��1¬�:��4�lm�:�f8����=<�>��.5!>�ht��G�2=Q?+ji�,:�!I58�� t�C5<M�wG@�@���V�a�6W\/\�����k��kE�5�.y��x�m�����=��Yg��kΗ@�	��y��q�k��PY<���X<E��x�
���ꉙ�)�!����[�e�������_4�i�G�p���T����NQ��F�\�3�`W$뇰&�ch�e<7�`~�/�W��U��ˍ�����+r�m�ˎ�=
��东Y^R0Wڄ�K���^�YX���M�w�w,Φox$��?��'����������m�3�쨤�#��<�	G�cW[�r�@�O	Fax6t�Ճ��A�B�'6	�ܰ) ��[ (8D��a���8����c�gМỷ'd��}*$����&Q!4G@��Ŏ��"
:�����C�K��^E69�Ԉ`�+h�Z�;!�}]�s�f,� 8��%�M�{q�ce��3����b49>S�g�C��D�����P^�l�X9~D��^OJ%+���L}(Va4
c��([�ϭ�    IDAT�!�߆ZZ�~M��C��_�5��-��>2y?�L����v�� oX ����� ����{�b"Xz3��a���?>i���&�!zm/F�ၙn�a��%~�[����a�Hm����-)+�����<��H�/	U>��ݫ|���@7~M�ks|�}a��@3P~l� ���`�l�����1�������V��=��{4�A�����-��i���>>'�1���:
ދ�x���hN�3x/z�C)AWɸ4��8_������jH:�������Jr�n����I.?%�l^Μ^V��yRj��w��� _�)#�䩃�v�{ǎ�o=A{Z�v������?�������}��K�1L>�.��P�
\ h��oX�c�aVb%70'M�,  ����7����M�4l��B�N& �M%h���d���~X%�;v*�PPA�?�4��	�E c[\XP �����K��no1��ݵ�3��]��(���@`��L�̮��gr����3_et�r�g�^�"�s����q=���}�L^�U	>����9,�R��0��5�L� 32LϠj���sӝ�c���*�x����a�.
ڃ��C~�H;�n���Z��Lx�y��- ��h0�Ԛ�\Bx��2�-�����H׼(8Cݎ�F��v��y����>�=��c
���2�Y	̕LBz�vk��5O7�y�ɚ��o�n�d�y{��K�{��>��+��f�Vk�w��Z��$����ϣ���X��:�!��VFsYi�n��iҦi�g�c�7oA���Z��F�J'b=�w��qFZG$����E9��$5��29������Zw�.��'o}��ZܔV�&�@�um����U���efz^zxYն$���x���?����ƞ]�ܿ�/�V��{���x����'��������[��3���3�� �"*�%S	�f-wbQ@���Q����AT  |�*`��+|��� XH���5a��0�0��בϬ9��:x��q��qk�R�VU �w0���ܧ�'t�>�`�c��𙠆��p=@� �.Mbd�~��QE�n�\�����	�>�(��i9��8�sxჀM�'sƹ8�S�\�r��׋A#o)��x8�[��]�n�@��Z,��*Ca*F��R�	������̼�y3�0��"n�v���a	����~N���t} ���i�ÀՃc�wW�}x�����Oh��1��#�F����ӌ����tQ�N��,?oQ~]?�d����6׀(�Zmp��a]��P��� �Q���`���K0GJ"���͢f`�{h�`�[���˱�ϡ��e4?�`��O�T&�jku,�B9׭V:+�07a�rCۘMOOj�1�  />t�aM�k���vX��=?7#�jA�)���wKqcY�V��C�el<������Ie��h���-�^�F�ڞBI$ݛea�(uݖx�Wݵk�������'��O����//���~���7���j��%�
�(�SM&T~CA2iA��A�,�I탍X � ZD�����}�[�����8`�Q�]�d�XZM����E��v�7,e
���/h��FU��2 =��
H/�˛)	Ȟ��̚���)^c�o}�z�Lk�1>�I�k�y����0���L{�1��i�f�ͪH��{k	�]��rY5s073�WB�=�8Ђ�ah6�5���470?�w(ʃ�}��@�B؍����X����?�����[��Ϸz����<���)y�3:�06�É~-)h����3 p׊
9Ä;Z���ͷ.����߷g�>y]B�G/XӪ���]����0�`;���Ѭ�a?!j��/���X?�«Z�B�*�5ӑ�Q�Yq,�Rn5�F"e
]m��!��7c4���#�c
�l�b<����I��z�4v��Y��kࣵjY�y�Œ�=�0�CN�:%w�W�v7.y��h�eaǜ��.�/Ɏ�	���_ZͲ��9-�27��5;��8.�fM�i��}��y��<w��6�q�������u����=�����뜁����_���憛n��F�#�tR�; ��� �uchJ��A�?��4�T�@� �́ϔH�U��s|b�5�>j�l��cǼ��	Ld^�.΅�]�tC��0NS�Bw/l�|PT��c�20�w_3���=��d��qy�*���9n�ez���b)�MxMǀ1�����a����9� �)�0�,`m�ms��2uk$���XQ��B���j�*WխE#�S��n��@BW��4��#٣ff�� t�����������A��z�u�Ǒ6�~=��E����G�H-�c�G��Y�h���v�D����	"J�i�e^ôl�<�|���!�{�㕱�f�< U�l��_4E5�I��0�L��Y`�����Vp�|�ɣ�u �n��ϱ��ݵSݍp�m	<��!6�9>3p��Eݷ��T�y���-��٭�{vfN67�r��R�5��`5��-9r���Ҫeb<-���$��Iq� �DZf����W7Ve}sM�zq�^Y_+)�7]�Y�i`G��xWh=;���.>��c�ؠ$�#����s�=T������7�z绚h�I��X������\K�����Z/�;�A@���
"A\���/��=�c�aR�f�� ��\\S;�5L��R���;4nY[ې�.�H��A�u�t�s��ia y��=��N����(���ϸ�7���g�^�i^�`eR���`M�$�qӔ�
���S�0�[T�����u3�%,�Y~���k#8� ֥R*�� s�,\1=_��|�`^x|�g��������!�Uz����r���(��g�
x������ڶ����GD��d��o'��;��7T���t����ˣ]�_Ã��G}� �r��ݧ��Q��4r�(�dF����k%Ӄ42�3;��\��o�zi����/WZ����� ��ё��|޽cA-���c�5�4^3�`���M��H�V�t�N[:$�\|�<��2==�f��o?*�RE$f�y\��K.���LL&�)y�5�)"����N��R�Wdu}Ū�-,J�P�j��j�7S<I(=�g?������(�~����3��O��_�ɝ�N\�B��LZ��QIg��k��R07��U16���2�l3�������} 
�`І�D����� 8CMc�Κét��{	���hp>�  8 ^4IG�=��j��f�d�g��'��k���j�Ѥ^{�*�����V����i��9R�3�Z��?M�g	a�Uc�8
�جK�l��
@]���A�|�������i����J�
���	-d	�Y�����s�o/@T=���agm'�i `��O������:�~��x��O����Q���P��#ωdl�-��G̃�ct�(�o�g����@�~�}���xh��ʡ��;��S&p�*I���`�j�J��Je{ΐ׍FE8�%�'v͇�f:�~
ip'j�hO�g���a?jIV�6XQ3���fvS�B�	��a�D���h���򢟽R��~�61>%��_��6%�A�,vٳo�<|�A4E�\F�w�U���%�+�R-�U(Ȍd�֬igJ����9�U�R*69�TS"�0���6�<7����<7;�X���z�9�OVw}��~�/�;~ꥰ�FRC��9���S���,��͘>E`���t�F_�	��`�@M|�6M�&U[kJ�
��������x/��V2BJ��ѐ!���t<����9~S�2���&ʨNFq(����2t~���qyS[��8nCs(#v�҇�W�9$F��Ga]��9i5�fn����A;/a���g]�d�cD;"��7���0��_�-���6w�0P��Ki h���D����2�{!����1'?�(�s3x0��iG������liL���9:G~|��]��3������-(-�=�@�)� p����5���rƞ�ͼmQ�/�,4s�9�����������TN*T�?�/���LOj��g�I�V�ְʋ s�HB�Ao��X�{�є��Iy�/R�&��P��z��7��53�1u��z-�����_'�y�%���$�ki�ϫf^kX�g$�i��jI{��k�f���*�����!ёtRn?���7��g�=�>x��~���O��O>��Z�~�y.��T:!阙�`bG��~;����?0u�F���І��q-�O���~H�<'(1��a�4�1����i�e���ıAɘLx.�G�q�
*�9S@ � �QS&�F����M[������A����[��E+�~<��%���k�Ӭ)�Q��@on�kh(���cZ���Q�`$�rE6�Y
"43���,u��׌Q��it~C{�� � ���0���ٝ�{�`��0�R5{��c�i���H�uTh���9y�f���07���Gӂ�	T�|/qo`,�p<L@`�a�v��Ef�~N�K \˖� N�m��<)�C�Q��fO@MB6�5����qK/CT8�bG��ZH½��� �se4c�x~tD�� �ˮc�Z8/ ^�C<�c��{���!ϽY��s_t䰜>}:u�����#o}llB�g$���'N����d�=y�+^.��RY_[��ڦ���2:6*�rA���BA��q�͒�3�.��<�w�蒦=k�?���7/.�o|������������<�����g8�|94�tn��=7�&v��@ ��{
�5�T5U��j9�x�O����E��mp�@� \��#8��=�>���յ�>h�7
�3�Z �C
���п<��P� Cf�+ީ���z�=��k;�!�N���̝@ݿ��/�vB����m�Nb�jS��Ph�
��{0@�m��WWW�q?.ZNu�W���VG���6]�H�T�"���R"�����4���}^�,x- d�8�O��S�
	}�2�1�k1����"|�	h��ͿI�"�q��L�����ڎ���g��Oa����_|��H'Q �����ati�^
��=�{��� J�56tì�'\�15jً��w�� ���<H�D�@\�*/�U�D<&~�847X!�j��x���j4�ȱ�V{ckW?�o�fO�Z?���)A�瑚��t���a�h	:'! nye�_^�����[y��CX�p
c}��+�N�T�k���J&=�9�/��j}H\��^��h��i��EW�+ᥪ�7�5��O�NK�R�f�*(�59�����m�.��!(_@�TJ�|�x���{���.�;��Gç����p�}�/������.���}0Ϧ��$�,͆�ɘV�M-�D�������|xW��zͼe�#j�f�էƅc�����?ab���z��%Rm��h�8@��lJ�T�`��@�X	���E�	��g���e�̯�Z	�9�������mlO�����4>�=Ӧ���?����J�.�5s�f���`����B� $p ����,LU�}rx�A;d=��@� �A2��0`&(���k��H�2� �s�&z�D�!e;a��w1E���0�-�̚ۍ��F���,DA��y�":O� �������qg���{
���{���S������Z���~�X�.�ͤ2z^"�W=�����MA�-KJ��0�X;���A}a=�b�T�SB��T�I��-�ۄi��պ)Z����}��hq���BK�zҪ7$;�����r��h���y5��7�{�n�hc:11%�JC��.9v��r��^��W�R������I���0_~�"�u���x,%ke�T���γF��r��cq�������|l�������s�߻��e�^���8qj�DJf�Y�07?���?�+�1�F�Z�2�CyhH*�q�qA� p3���&&c\�4C/��\룲q,�)cۿ���������4yMfv��X��#�X�&b��7��I�M���z??�>?^|�A�$�d��1d(d~�/%�R�pfxsiTK����x}>����>!	���LW#��d�ԆX�Zg?��f);V--.�P�o:ߑ@A���f��A0�'��V3P�\yaJ������5����	��לs�9�N��q�H;��蹏��<PШP��4H!՞��
n�ݻ�<0{��kc d�����M �uT�E� ��7~-�'�<t�q.���1�!�!����8������5-���f�A'���,�SԕM�	��ْA
}� �;�N�V�u~B�+��o�>s�� �x����Bl�b��Uvț2�։P�*ӢY��/�\V�#�{�.(:�g�\�����s�r�-��=w�X���}׼S��s���̤���D!�5��T*�>�r�����2ӄ󠙇
�j��db2���d���ԷgGF���"�?��9�o_w��|�s�����#`��,66�Ӻ����3�g�� V0u�#�I��4���G��G�% )��ZH`+�{�	07?��f�RM|yY�U�l ��U�Ë~p�d��U��Q4fϞ=*}�)͒�D�3A���"1�&�i�ܘ�p\;��p�<� 4+�zs&�g��8��9�x���c���`���̮y��Y�rXX��x�>0�4����u	zfF���{�h�2v͘@IW���k����K��^h�x���L����<�&��X����!׏s�ז��{y͚���G5_~̛id޲��5L��NȈv�%�<�i2�\�6S��4��~���f����L��t���H?r�?H~����n�0���ʃ놮-����q�����;5
�e� ���!�DR]�b�t F���+8�L�1�fv܋��l�l��^��<��*t��ŵ��LV�˽�:�&S��5��ٔ�������#��3��L݋P��9>���aL�(Y,�$��i
�]?�U�����}@Ӆ˅��gT�Dy�J��Y+��F�eu� �r�,0�Z�}�+�nS�Y����J��e2�e3�;ڝ��d"�l��I�I@b5x���X)��:�d+��u;�^+�I���^���v��i��RG���$"��O���Y�朁�׿������g��A��锚_Tc����~���ba�V+~��fZnP�.1cc�2��΅~��i�ӓ1�����q+~B��=�B��\�����J$Z��j�٭�LO�Fq>�}��19r�n��
܇�;�����(�"�����ҤB9׳4C�/}��xJ���d��L��*=0�yQ+����i�����̥����n.���^��}�^���|^��
M�����2�L�O�2G~  *qڝ�h��G4�`�\�(���(w	kA�l�ܯA��O!���\�DtL8_��M�q�h`��a���[�Q�����I{����HQ:�t����[�&�`����0�EA�{L�Εm��hY�PO��M��p};oP���%(@a��Ӥ_koj�������c�f�ǵ��UE<NN{�f��ښom.'���Y�x�cˤL����yvdT�G���������B����*ժoֵ���{���ϔIk��|>'�E�����$�R�W��'����{��dӲ|zY���)t������Ȩj�+˛R,մh���Ы��fvq��[b�ڪ���Y�t���X���Z�x���۽x���{�^+ދw����%�����8�k�dr5!�r,/$�j"�ڌ%c��X|C�[����^�[��2�TK�҈�b��x�_�̿�w7��o��[��Q9���fd$��E�A3Ǆc���M ������W��B m��6?�6w�
��֪��82Z';���
o&������\�:�A, VX 0�fv���B �݂�LR�yym�kRq��7�G�,����L�Q��kG<�).[����~�F��ʆ������7� s[�V���,2f����̉s�kb|\7?c& ���L3�e�y0	����K�    IDAT5/(��8���� ��u��[����*t����an���r��q
[���D���G!��*��q�vP
y  ��HoK1'���1v���dO��i�Z&������_�a\O�;�&9�`gfks��̎ߩ1�^16�T  �R'_j6-u���( �w])�G�z�=i�t4<�9�,;��2���1n��t�b�-��\���� ��'Ƣ1-m�x>��F<��i	���8�i�_�͎s(� El��r�%�Ν��\jvOX 1�N�KG�(�Ӓ�w��e�PTK�-?���<~L���7ʎ�9Y:�����K�Dm�$���jޟ��냹��u�B�i�8kܳ��XW��&�����l�
C@t�l����sP$�����X����d���u�x��J%V���}�L��H:��L<u��L̪�=�s������_���Q(7�!Ս�G�fv]�`�q��-����)���A(ls�y�f�DM]|�XᏥ�h�o�8 V3#�Z����tc�bj�Q�޽G��ؽ��� ����ܖ@x �"���?67w�F׌��M!�3�a�\�"�\��Ȍ�8B� j�c�gNZ�CO����`�'As�\�9��GP��s�����L�T.��-�9�1���Q�8B����
�����^�����#�k��I�:������k	̂2��t�NX�sE��?�����ߛ�%A_} {��w��}�`��G� B&������&cjd<��ZKz��:l.자��9����G��Ҥ�� �$J�>��y>���`I�T<�es�8�%�o�~�F�$���A��>��"��\3|���Z��aMP��cɦ���`\&�u5e�_(0���afW�(���ֹ>k�̵�)�}�A@1ƟNZл)#�~����c����׹��U�Q��z�s����R���̔\�^��$*�5���y�T�:�ё�Z4�)�����^SN<pLN�<.�t�/j���3�*lLN��߽�*��ʒZrfgv��Ҧl���R������H	h�����N��ۺ�Y���]�k���%�>����w?�� >�h؄G�1����dN��$��s6�񩩑���D>�30�� ;@Ŀ��k_��w��\�NB�ˏ崜+@Vs�C@M�Ԡ@l`�܌ gh�&�&T:�#:�����M�hZ=n#�EfK_ҀI��ɚ�n8ǴB��--PA��;֗nq���a��č��Q��~oJ���S�"��
�Mύ�ϼP�5A=HF�+���{X��n��X=qz��N0�̖�4�������4g�:�:�I��Ҳ
�e��0�{��a~l�� (����ٳz�����oߞ�xbei�����C�Ri�^o�Tj�q�Շ�O��E�3 H��nO-=hM�t��NեAa@��N�{A�����^��ԙ� �9�5䩑R���5�?�9�k� ������� 4�l\sާ/d v�Z*�K{�kG+�d�Q�Q�1/k݊w�g0�s)���;���gj��t���.�w%�ؠƒZׂ����q/�TV�	�=�O���t��>���sj���Bs�f�S
���"�^0W}��Du�����O��JM5s��bCp_�8t$Oh&\3��l�r�a0_]]�ﰏ�U!���p���|0��޸�"�)fx��i(8	uGb�)�g�9S��V�IiN]�+���B�(��ϓRiC*�u)�/�կz�ط[J�2����@���%���܂�.�iy�Fа�.��	�fN+��t�s ~�1h����i\E� ��>5�a�qz�HL�]הP�'�9�]�#��l��5������X,�3���9�����O?���^��7��b�=���t�ɤ\7c`���3HG�H &�zp�3Ԩ5�<��*e���C�$3���7��	�aL�1�����Yua�錿SKŸ��+I�<.�4f10����	�Rܓ��Ma��l���������s_������.����.��j	!�&�`���@`���Ш^���b빵�6'�f�H����kG����|��~��?�`��w�������c��ՙ�����r�����g����ju�R�̔K�I0�z�av�+3��Ϥhl>A]C�2,��D�Kܹ��3'��|p��uP4�ڷ����#��{�����#��2�T�?{_p)w�.ZbR�ECL�.V��@( �"'�P!}
�Bu.�*YZ 4ߖ2w���Z�
�	Z�k_��)���P
ή���϶Z� ��L3Hme��xhQ��Y��0�Y�0.�E��^�&��G�'�
(t�p_�}G�
4c��41�e�i�&�cu1~v]����ݖYY���U��I~Ĳv�/���J1K#C�8��fP��(SS�*Ș�����y|���ƿr9}nt��ƌyT�)�R�Tq	�Gs��\O�%�˪��ɦ5Z���>G�/�bq(Ɍ:�ܨ�k\MJ�ݒ��eW��ϹT�Ϝ��/S�S�,"�
<��Ս)l���-��������+��^�ȕ���b�r�G�$���y�U������!P�%ٽk����}��B��'���O�z#_��W��u����j�n"=��se�b��٩	x����!��`��-5�"�?����zPX��2A��Z�o�����{�������p��C)ۨ�Ka�kS^���W�NfA-���櫋J�L�"� @����33�56^��63�U�+��j�C�v0+0K$sd0O'E.����W��{���|檫X�y�5`v��;&VWK3�B�R�xhm���J�t��J�b�<_(�R&�X ���5Xq��4��ȭ`4Q�˴�A�?>s��P��
~S���6?2^h�}�l-�ؑ~���DiQu�pn�t��kU6�  Ѓ�N(4� #����}&��@�;{tc�)�Q"�����;��@�w���i*�V
����R�TP�g1M��z��y+�kc�@@���"���(�<��L-[ˎ�Zj��59V�M,�R #`p�P�H5Z�
EU��{QР�ߣL* �E�*�=7Z���"��и(&m�0�	�J�'|rjJ����A.���Դj�Z����<��K������^C��C�KgӒJ�4�/��a�:��N�Gd�ҙu��-R�_�<����R6V��L��䌌�'T��
r����7���Y(J��z0���źrmh��5q����*y�'�ĿE�(��C+�����2?7�Ў]�o;�s����x�;'���zo�S�~��pí�ި� ̱���CR���i`��P)'����I�f��'Ҵ�(��d�)����;�DtI4{�w��	��@CA�hy�>S�0P��w��o�
��v��e!�3z���GH�
�! �_��a�a�������	�<�sF�9J�j�n��2K���U%D�s���Iy�����^���xի^p�c%��o>6���������յ�+O=�t����b�R��I��v��F�*�tLȂ��k�뇒�!��~�
��y�̲`f�6Ln��kB��߮2����t�X���fC?W`�,�.'���Ia+�4
�����@}Z� �?,`pq XWtF`�x)��Ӝ̘��0�]��7'C ��e(07�������y�{Z���L������}���p��.�R�kje5�H�3����2���6��A���@��
MXcq}~ ]qj1�u-R�i�Α������V`���=)���M�Wjr��'_��W�X�H<�Q��]�lGt63����t]d�0�@,�C3�f�.�t\:���R1�$�"B�"�Z�`�Ogs��|Z��M�v�r�E���W�\*����2�i�]}vľ��Q��|sQ��#ed������@�}���F�|���9��uۊa�)�Qh�w�jQ��ƪ���<|`�/+���s�g�1�گ��n��3���=;H��fn/�� j�3}��̬�_<x|��#��Od\5 ���L/���m�I���#C���&�����/�g�<��ΡV@͖ �w�`̯���!�
�J�.d^�5�7K����f�Ѕ&�a`N͂��3*
�&�a`n�� ��K0���˕W^�ɷ��u���_�:#�t�ݳ��K�++����>s}}�͍�b�V�.���vw��n���4���x�	�<�w�੍��	��ܗNYV��.|ρIO\W���}�ƀ��)q��(�aLF���I����L����烹���9$�X%2D��9iރ$~�V,j�L=���p���sp\S[��B�Oˍ��O��`ֆ&��  �s&�m2�����8�a�j���bp.*�yA��8*�W�+��5<N ,���-������2�ׁ���@�I�5/XC��I��[���d��hV�Q�H:W �eϔT&)�_�}y�K��뮻^n��6I��%?>�`n�k`^\�SA�\`u�5[ '�NSF2Y��.Kg3jAA����V�p����\C��A�V6%&ٹ8+�y�+�ZF�`K�1�Q�EL㥚L���5�B}�����,Ѕf�����a�D�=�$F��_�,hg�9��SS9Y�9�.:4�/b��(��뜀����v��_���w��s��A��
w�5d",�f2+�Yt昴�5�����e�F�	�����/���ظ��&�DǱz������q����Эldl�������nA:��*�غ�\G4�N|f��#K{��C�s��hf�6�f A�ͷ1�O����z���{����;r䈥<��ɓ'G�_�\_ߜ*V��676����
�¾B�2W���k��h�^ϷZ�\��Nt;f��w����� I��#��1̶�vƹ�Z@�Kj���!�p��b����m�$�ʁ��<��u�/�{�/4����h5�r�֏�S��i�d=p��~3ߩ:�{<(�2�/>313H�
f�|��[���,�E�7�U�}����s�<˒Ѵ�Y�>���8���<�YM}�Z�
�'Й�݂s�z|�|�|����J�Z1Ҧ�"5�v
<p��r|�2��'�FEV��d|bT^��K�Q�=������^�������@����R��dl|Jv.��1Y so��}�L4&��J�U��HN}����a|t\ߡ�ï���4��Qm� ��
�8��mI�V���	y�^+�jE�t`��1��0N	A��k�
�'�9� �1����6��߹o�/�;�V(=_��J�B�#N�X,����W�..�{|<��$X׹	���3�?���|��N^�n%$��k��/>s�E�y��D�w�`4?�~Q�bB���@�����9��{�Zt��1S�!���1���$���b�qs|\@��_x~TK�9^`��=}�d�[����xIHQ5�N��&bB5$τ�#th&^����g�fZ3��s�����Y"J[|ZC�<��Ɏ���+^y���?�C��,��)~;vl|e�2�^)��6��Zig�X�۬7��m��Z3�Ry�RoL4��	h��1KPO�o�(�ӌm�qI0e���U�;v�Ai���[m�����~�Z܇kAS&փV��4[Qa��B׆E���c`���>�r̴+�	��RX�|��8��F����g�3X�TQ�I���շ�1��}m?&U�V �&��p�l�@��?9>� 	�*�8Y��τ}�s
8�`և��V3
��:�����
4�"Hk#������9�y����mxdh�9V����YϸTv,��ާ y�5�;���\q�r�ͷ�3.{��z�m�����l��2���;��9�zӄ�(狊��0~�mͤ t�$�(�\N`iMAc�y8ד܈�� ��L�����rٌ4�������oz�4�5IgR��ZZ��H~u;������̇m{�9��R�J� �{ߢ�lIm���x��KK̆@N�C*: �����1��}��05{R)j�D3���Ǐ|���N�yv��<�u��\X���/���h!c�����C�X) x0�B�A��̅`������:���K�K34�A�`���;7�I���.U�̜�L-�ob
�O�/�f�nY<��`����Q˄x� ��"����Z��&�?tL3�7�gn�?%�DWf�6_s�+~�c�����c�#^�رc��v;�\mMT�թbqs�f���Z._P*W.(����(L���F���F`f^�G	*K�r�5!�s�s�iL��щ�1]c�	�%fI�8���A��`)=��m�OZ� ���u�q��2ȑ ���_I�ⱸ5s�5�^��h*�R��1��d�^�k�jnN���eII�v��ι���f������ p3]��V��Ü1�1#x��5�?�R8A��6m
���J���P���y0�������x����	��٨˳/�Dr#)Y_]�N�.�|��4����/�;��!ӳ3������?�CKEI�����\l��s�֓�<+@1�L(���3/�l\S��w,���l� &�m�[�RXL���Ns���MOf%�B1������V-*�#F ��H�c��Z�R�p�����a��ꆍ�s��Ĭx�#�+���f�~��wh��u���B�A���$d���{��}��L�'���	���'�?��D���K�Hu��3OgL+��<CU&���B&'�ꦋTO#c�� ���`g��`����>HC�����?�� e�1RJ�V_v�'
���N|�-�2�j�	��	4U���� 8�+�[5
,(l�qMJ�f{Q��B��ϼS�h�@ ���,�}��#&���S� ��۵���W��w>��w���OŹ�^/v������ՇN�ll�.��>�X(\�����T������z�9�X-~�|G8�7��qD�s	��d�>�ǵ2 �S?���ݭRI���i���,X0{���3�4���&i��H���,��S�ц��Z�7��hZ�0�u�Ӈ�68Ǫ2�(Q8�$ ���w���t��L�j<p-9���F�|&��:{4����x�4J�k�� 睚�v�V.�k��r"�����\Wff�J:���|��r����'Go�͍ey�5o����er*/k�,+��������'�ԈLNL�e�v s�,=c���`�Nu�}�{���~�a����ha�d����'2� �����R���S��~�6��_�r�� ����5��V�z�!���>�$����2�<�|����|9����1��
�?s1W�<���XGv�?����fg�7<>tN��~x�_������C+Gⱌ���In4�f��㒊#����eO�@:����I$(�RK�$qs���f�7O{�Ӥ13�]���@��l`�$2B�׃:��C]$j������d�d�$:���5B�vjF~<��>��8wl�e(X��ڱ{���Ϝ��`�w���`AA��`�J�UK�a� ���LZ���w,�X[��Z\z�_��?�o�������n�m�R�M�>}fauu�`�X��X�)W�;k��d�Z�wڝ\���tz#�n7feshI����HD�c�#�������UXS�Z�S0�Q��4�Ȩt���;�
� mI+���co)o(�C���o8���bM��q����PF�S��qDõ�AS�Ǿfef$��n4��
�Z��q���s4^� (ۯ�0�8��>16Z.��Iø��q�4uv/�s�hv���`a�s{]=���B��3��;��3ט�k�Q�g^��LV^���el$%?��u��������r��4�%�p^�X�k��e��o\'���&�m��0����Chְ��-�L�啯|��띯���LNZ-haj��=zJ���~=�3���=�LN5�v�!��K�V���/{�L��i��<jI@Śon��;~k��ꦔ���5Ä��kOeC�%/����G�ۃ=�0�/Ͽ9����\?(D��ٹkni���w�Z�~���s�����������3˥��nRr������J(# �I�]��Ai�>0���̂�N%S��o�=�    IDAT0�����\�0#�4"~��Y2.[,��A21���5��"y���r^�3بԮĕ0�׮y.M�d#�`�����`���?f��af�|�hy�׻�=}�H�;��*�D����=�J��j*,J�:r���Sox�k~�W����l��^�B{���&67��Z�0^�Tg*��|�X�Y�Twժ���jk�VoL�Z��N�;�h4��z[A�wļ[cT`Km)�ec/T��� � �������Rx�<P��*u�Di�*����p����i-�8H����4��G���ܫМ���i�t���H����ղ�R�@Lc�s�w�V�9�@����S�Ho��Wh5���S�ýM3�Ыq�J�9��0��P�oΫw�l٧�?�kj݃Z�_����*|3;�ᅹ)�&et$)�Ҧ|��&�{��;�j��ߖ�W��7�&_����1��c4;R��9-V�mX���z�vE^���G?���
i�[V�N�t>��i�_���ni��X"��bU k���}�d��)��%?+���b;=�v�V%f77�Z=n���(���aQ>J���4ϗx�c�(��:D���a�\�9Wص8��=�rO���0��|��������F��3{.?�`���s���7�5??a
�!M%:锌i��y&��h&)��=��2�S(5y�KnQ�ٛ�	�ޏ��M?�ޱQ��yP�Cs=-�A͜��f}2i}ΐ���h��ٓ�M h5~s�lj��}�?hV��E���"�>?h���z0�f���6�>ӌ���=�N������;�y��{��mgΌ�Ry�Ri��JřJ�������z��R���X.�֫��F�9�nvr����!#�td���u l[)R�gMS1�6:T)�u�v�u]��}��C����dF�����԰q/h{x�
����p:~��W��A����p�9,u���㩌E)����Z�Y�,���� >���a�\�NGS,�3@#���]�*a���w��S�����Ѩ	kP*�M8|�1~ �P�sBȅfN��{	�+ת296.�JE;���Fd��y�/K&�3�Oʛ��Fyɋ_,?���e}}S.��r�=��G���~|��b skT0W�:��`�#0��_嵽���M�/�쪾	�����O�m}~t\ݭ�nB�R_J�]��G�jyS굲������ࠖy]���\��+J��k�'!X�)�˰x���->�_��AOtmp�+�G�M�5s/�{�5� H�m
OG���,�i��1�[�M��O���0�Ե_��o�G�_.wfzݔ6Yɏe�!�k��mZxW���$*�7}S� ��_��4�! %jB�(��9� %jn����{0��@���Q����u��OF���� F/8x\�"	����Ԍi���m�4ا�M���<�3��~L�n�ܪ+�����"�z}iȍ��Gs<���d>S�����y��o~�G���W}��l��Q�=~�x��Ύ
��Rqn}��gsc�����%�JeO�ٜm��3�f����	>v5�f���X��fG�G�h@��Zs� �`�1��	�Xc����׶� �R�0�_�/ߛ�q-�-��
���ƹHe����ڬz�{��PzO�m�	$����:�����Cn<+�E�YSj�i��V"-�<*����Uc�q�3!u��N���af�L�)�z�\��`�Zĥj���l
���m�\��l:%���/��͍UY_=#/��E����ѣR.���K�!K����"G��P�5, sq*p��c^����7
;�K�����T����nd�T��Jj�o�1,����4�~�DX�T"L�vk�-�VM^������Y]>%��=kJ�Œ��]_+I����YYZِ�BI���J� ���m�U�<���n; W~�y<��Ac%*��s�\���Iٽc��<8�/�LF�S�^/��O~�7�����^���ǲ}0���J�!���A<h��YΕ�+M��ɦ�l���ƨE�n ��H [D�������p����4eF�����E�1����a�	h^3� ��1�o14� �����V����p��7���� ̣D���	�����;j�07i�M�fM����nL�4����{�;��o|�+��?* ?��:z��n���|z�ܨ(*V����|�^��j�\���J/�m��X�{�X��Jz��rV���2�Mi�����K�������K�eC���$�FZ�:4I���Pv`�o�f��2I0����@_oT����>���y'j W7D�����Z����FW���3�u�f6gi��YSY��5�w��M�Ž��U����7�m�R7A
����h4ͅ�Z�Z� ֓�.<"�y֥��tJ��O���^:q�4�-9|�"�Ujr��{����\!tX]u�MC{6�i���șU�뗱yΤ�j��3� (P-�h�ˋ6iIk%PtS�9E�@O��"�fM
�Kr���k_�r)n.ɞ]��$�R�H�0/K�ٓٙYY+��꺴B�eϛ��pi顀��(�x|������Z�"SSc�8?�__0�ϞL���Q����W���G?V����䨂9��0��̪j���R_Jr�g���`$#2	" ��s��m3Y�L�7�g���������=y=l,�s�ySC�w�d40�z��O#�C�?VO���9^�̩ٟ-(�0�{A����I�~#�w�3���6>	`3;�2L3'�<��_��-~�k^���4�N׃�����J�f�;R*�Ǫ��l�\�m7�s�Fkw��^�Z��fs���u��|�V��z�R����-�����4zW5�T�j-4�<s�M����A�
���*ΜOZ�8 �ޏ?����T�O�U� -��k)m���M�Z|$f�24�"I���cS�?t�[�&qh� �4pE
J<��J�Mi0>T0�/Z�( D���&��������¥&�U�C�S�iwQ��!��'Sc�A|BR
Z=������5 nu�(�ł��(��s�~� ԏ�X��v�bA����P�,�m[ryd&b^�W0O[e<��h�D�`JZͪ�:)����{�����ь&ѓT:�)��JC6֪ҨwejzA6
5����VOK��,CK��+o�𨢧�F����6(~�5s*) ���,�N|i����LN�6�(�y��|e�7���}�_�|�=)W;�t*�`�hv�9
}h{ �aݹ�����櫨���t�
B�� �^�7)̴i0%��{X��Ӝ��J������0�ix��ҹ_@2jOԺ���lB�`�	�L���9[��G�9	�D��=��K�9jSc�����ԏe!
fv�[���S8�p��'�]9|��;�����+^�o?�M�O�<4�����\�Q�VK�r�=U�Vf[��l�V�o�;��U�U���T���w:ݑN���©-���z�V����&@
�V��(0,=P��a��"ﶢfNA��CA\�2����F���5s'-z��`�2
�������])Y����V�kA�H���)L�.�����½�������MA�ֳ����"N����7�q�F�p���g��i�ڵsAFF2r��R*原�������;wK��Ե[�,����{㟡j^�HM3!�����U/Ҫx f�?��0��])a�Z��˒�P��K'�������5���Td��|���Ҏ�)t&DC#)���V������J�)�YQK���G��
��
И"⭮�k���;�{� 8+�n0K��[棣Y����w�cn4��JR�`���ܜ��_|���{>X�t$�A]���U���nNt�@��N藍��#�3�� (�G����I~����(��S������;?��,�H�� ;L��Z)A���{R˦�@b!X{Mă+�c�K���
���%S/��W>L������j=�>�8f��*�1�)H�^� iy��cD����}�fι'�5�^�|���\z��ۮy�;>�җ^񽧘��s9��������OlV7����x�^�n4Z�]��u:��v�5Y����7�m�+��L�0s.�,�@F����ܠ;�����|��OI�R�r���G>5�aM�
f�3��A3��7O��j�)�#��h�јł�ȴ�^ ?��������Y��L��֤�W���\^M��B70 r�Cxa4
�!mI��n1�MF4H1 �Ow��)cc�r�Ňum���<nT���z(�JRm�����B�� �#��ܖ8�g^��כ�R���g�Z] �A�c^��{�F{kxWL�x�2�OK�U��Ѹ�������U	e�%��(j�3G��|~F�͎�>�*��	Q���������v��h�i�����j�,�\ZfgǾp��ON�,��	��r0�����>��?:z��Wj�|)����Q��E��3���P�/DA"������ $J��@��-�����Ҩ�elbR�Xk�}fPoե^�鶪�c�|(Bӓj�b����Di���� Z�Hb���/�<�{a���H�Em����E�_h
6^ X�;J�^��}yo2C��Qa�k�M}��㞼�jW��F��;�;M��xs1}S�6ץ�H��i��`�y�ݵX+Ls����S �>�k~�y/|֍O��z�c����Ӓn4V�<u�Y��{��?�ڵ�B���e����T S��a~�&>���4��7M��UL��k����0�ǀ�I
¨)�T��S	I�CkԎE��|�r�2�-�F�WԺ ����	ޝ�Ɓ�e�����#ꑧ̂�}Ƽl_LA����ĥ\�h�>|� 9Mm��V���+2�k��j�`�ZݶP�LdnvVv�Z�g�FM���O�g�|tue]A�7d��^�
M� ��|�g����+enn����ZV�n�ǡ�_�T�t*�{5`�GD}�c��䋹�ͥ$�A��|���];'�].��ĝ�<���4ZmI�3�J���C�RS�����ʋѥ�p� KK��Z�g��趈
}ˣ3��\���k��r��s�R�;�nۻs�]�?�-9���̏/���g��_�����zSFr֤ A��4r͡e�t�.<���rh``>0l����A4����}�ᇬla�Z�-��Y�DR���4	-Iiǁ4�rtD�w��*,���>�
E �� șZcR�����ŵ�j�g7���HA�7�Nl-���y�R�ޔD�!��"y�|���ì�.��chY C�oQk��Aj��p���N���m���j���	��T"n��� چ�C�N�V��dB�q����������[��&��y�o����_r�w����x��.�<�O-�sFtt�w@��;�X��hT��a�2`����OFq�%�u��G���B�O�O�ݴ�C���Ӄϼ�mdc���2h�S��߀i �-X�7z
R��g�V+@Ҫ�yK�����j_� L��.
�84��<z���.�5��e���cc277'�yγtqb��w��J�����D��Ɵ)H1�����Fh��3"Ws;6:���3V�@�5ٵ����"�<c��#9}.��Ϗ��X~Db��$�Uy�{�,�-H2ދ�k��Ⲽ\�r��BF�Օ��Ԫ��x1{��Yr�Z�b0WsZC�� *\Q����}�Q0�稕Ճ�6��d��Խ���޻g~��n��������w�g�����w�P0��*�B3��g�� ��2�`rK�B3�Pli�2r �)# ��7�P���s�X ���O&U]Z:�D�sqQ�[Y:�D�G:���ڸ'6����;v_��K|~Q���Ši0*�^���D]\J~^�؎�x.	�p2+/Y��6͐���y����)������:���گ�V��c} ��W�Q������H�����g������|��/��n�����f�ر��o��÷�v�?��LB�f��O�8���M�>p���� 혌t:�o��`��;\u�5�Q�ɘ �-�����
�b��w���ʟ��S�$l���ުD��wTp�{��y>\Z�����ֻd���x�!���4�`���P��Ƃ%L�z�
���;����|^���*�������>x'�ǜ8���m4-M�����GǘY�P6�n�
^���,��|.���̌�� �lnT�6��	��̬
��ɸ�sy���Nv%!Uy�;��K.�+	i��Gz)�&��Y�������YY�I�l.[�-�*?�Z�w�sh�S�#���ϟ���c�,���F:�0?yfq��o�ۙ{��2�r0��|�s_��O�~	$������4� �*�PJ2Hr��"+6�~0�Ф�Ʉ��ݐ�=�~��@�������c�`k*,���fo�,�g���E�p�OoǎJ���-���D���s��u}��ć�/(�{F�CߝQ�,(iG��|�����#M�ԼU � 3�sC��3\�i������c)W0i�� 7��]�XսD�)0ؔ(��g�^v��������\���S��~z4f��_��5���M���n=���SR���+���Y@,CJ���J�t�;����!P5���V��$��*h�fv���g�44<A3Wz�Y@hL�~%$Tn����8޳�Uk.Cp�� (tr�0΅{�[۔�iZ�ѷ�N�y�{!(/� ��*,�s�GH�R�7+���nO2��,..�޽{����i����.sm�b���-V�`I�fnq
!�!�?�_uC���Д5�/D�'B<-��)�֏��q���9ٻo��{�:��tV��r2:�5��^��r��Η^�n=�{)5殮���Ҳ,,�N/.�NmH�l��z:�:�����B
a�o���a`>l�G��ɷ�z?�f|@�����ڎŹ���yc�F�?F������:���|��N=��&��c�3ͼP_�S(2 ��4�`�F, �9 <�R!�x6?�:�h!i��a&�V��j�)W8��[�:tH{@�l3>�Up.MW���z_Ӧ��aPz���i9����?���& �y�����rO�v�=�z��vm>'��g�[�ڻ�,x�o26
M>X�Xؔz�j�3�	��B�ؔ�e�z��%�g]p�{�m�첋�>F���aO��x��g}�������s�,�jt44h8��������Uu]����7Usoa[f
*H�o�baMs�=ڃ��B�zM�©�����֡����Y���X)h{�Mf(\�������6ܓ{�&w
�^X�~B�q�� >v�c�6 4�~�С�����<������C1����Z��
��7��M5��0�+�E��W�1[&�
��"
�ƌ��R�x&�FT���� (Wk��(���p���/˫+:������x>-�xS^�ϗ+_p�ĺ��a�cc��Z��O��;%���N`n�����-[̉+�R�z�w�k�Qa��ԿG��/���P�y$��"D���(5<?7%s�|ၙߊ�b�'�E�r0����.������K��n�� A^2i��{��M�Ӏ0�Q�� F�� �TJ5p0����~�$Z
8p�A:�� 0�䇲�f3!��$ѵm�n�d�B�jK;� �D��n�LF}�D���gn"�7|��'C���=
��@��	Q��vDG��<�Ӧ=��x��/l�a���L�d)`��W
�~[Ǿ96�V8����g�- � @���}��{�w���w|���\p�� ?=���-��w��?�����^�Y�*󇩷�Bp�1r�#�H����O�1���Fp�5ˀ���AvK\�y�F��Y?u�MZ����!��~ڹ��
�o�j�uT'�;�{��i� H�6 ��Oc�f�'#��G��ZxN+��@@�n��V���|���s���Q��bN�;����D q_! ��AS�
b�^z��u���I�R�l.���&G��XO�1u,X��W3����x�C`��B9J��݁X�h��|�;vL3�9?>j��dq����^"����I*nUBQ�;O��FMx蔚�
b2�    IDATGF�����?'�SAav��ڭ:0gE�(��[�������������`�$_�w�Ҧ��N����_��0��'�k���������k���?_]+^���$���b�g�(N�I�S����{@�y]���^�Wf z��H��4Ulɲ��r���Ď��=�؉�؉�,�ĉ���ͪ&e������� Q�L������o���{p5�j$[ʌ5�{�r�󟳿]�m6���W�+�p���*nt;����h� �	�+���L�u���]�ȱ�X����I����. ����h���5o4��Am����o���J���/�@{���n;{���Sh� ��W,'	n5����hm�b��$��>��x�����|�3`�w�Lf��
�AM.,p���&$ �BQ��C$T��&��ѽ۾�?�������s/���z)3p�ҥ�G?~��S?��������"���E���kDH�;XC(C!(�kp1�5.ʿ� �9�H����Yq�Ϻv���^ "#C#o�� �Ym�i	`ԇ��W�ݔ���	2�(�FTro��Tj?�)#�r�J��w�8>䠙/��	ڐa���(V�,��������F�6��t�Qk�@S�27��
B(������(!�wd�\��Mu��qODU��;_�2V��`<������M��t�,߃����C]�aX�%9rd���u������v	�x��Nez~A=
�HB�fR�˂��	���a�1��ii�á�8}���m�ٺ/l�����ϵ��v`�q"�������W��Pk>�R�䚃�W�r������w-.e�"��9-s$<!1�2��.8�)3��M�X�X\���Ub��Y*���.24���B�E�[��
+<ͦ��� �R6\��@���H
��b�~�0[��#��l��vqss3��nAjh�/��O�^����)XL�-�����*����о^��j���0�7������q����xG�̿�-�#o����ݡy�C�]*u�Ƽ����������#��$�ɱ�����z믍���R6��9/}�������G���Ӌ[5��5F�u����j�w�x�v6�';�9׎T� ����U�rh�@< P@���; �6mQ%ɒ���>8�k�<�jy;�]ݏ�h�Yo�k��
H�Y��c���9�d��^���G���{@K���X�&��8>����NyZ.gJbqm�9C��V��$���W�(�� %�<��RE�I:�K����Y恰�Q�OOJ�pR2S� �C��ut�����P�`,�����^��H�i?�k�;<(�{�.��-��oz�x�(�#�[IcRٜ����m21�(��0G��=�m�
�a<�ܖ��qE�e����[��o樢 �ugGB::�On�{{"�2�����`���<��O�����dKC�_�% 4}Z��U0׍�Q#e6"��������0mjh�j"�nS&����]��.�Me,~�^�I:P4�����s^Q�@��}�A���[?#ȷZ�|.i��� j[¼]I�;q�Y����"E����L�ak�������}QS���k�㱭|���y�?�i�
�RQrEt�2ݶ�6m���y�
�N����_ҙe���RN�H�+7����~ۛ~}̯s���<����gN��Չ������f�~�WW&1 {ð~A��5�J+�p��=��V�c���}�`k��am�s|�w�^ڨ�_�,Ԍg�k��ս�ʅ!58�u�L�3->M8 �im�@�(�H��KX�y���	��o�}@�È��I&:�e_Q�R��A�
hQ)qmX��^�P&7;<��y�X. �,�(]��VÄ���̹���Q��p������B�H&��a��Y�SSS�YE���Ԕ~���ds�%'q��+�sG�����H6��Qh`-�E��ճ�etT&��23=�1�*7�#ɒV3~�f4<�4ւ�g5�M��o�aXW�s[�k�*�8�A�^�����z��EO��%U�9���������g�l�qX�sd��;�s��a��2$x�"R갊�2���3��f�f�Q@`aT ]�`���6��l�g�)K�" ������/�USk],�լ��a��l|�r��ڌ��"�+�@L%���� Z�͒�f<��
�����®��bBY�I��S �zIFb2�e��yǏ��%r��y��׾�ޚH<�	M�d\nؿ�����c��eˆ���~Ǜv��Ug��'N������i9�?���6䲅�l.��
��%��A�	��!Oq���R�dm���viI�i���4���`��T��w�.�IM�b�ب؆U��Z���Lb� �'@Ry ��; �&K��A@'Pq(@zL�[��
��
��MOo�ck<�$�`y:ml�ؠ�7:аO}�T^IU���d�;��ZCJB��e�O��34�f5�Q.ZZ�:������2��6sxJ�0���k�v�mr��U�d��d9����z<eJ���z�$�nq�@n���.������%�2�U�s29=��K�[g6;)[�H�j�9�#։��^�[�7��l��n���osxO�Ҩ����sl����z{C_~)�f�����ʿ�����\��@�`,s������2$��l8��fRH8�����̂4���
��.5Rh�
fN�$\��:͸�r�ul6�)��5Z�L4��h}�/�C�H>�ĭ��A]�Ά2gS�9� m����k�~�RD+�ϥ����ƴp�bnu#�zl����C`�RK;T^-s�O$1i�%d������n�X  ����/|A&&��0(�HP6�y����������_�X?gmf�̙�X�[N�R��La�;�\ؘ�dv���m��T��b*���/-�C�l6R,� �X4a,d$����dB�j�}�J����ڥ+�����=�0�>��iu�5����*��H(C]5�E $jY�n���p�"��>rmBkWVZ,��ݎ�lb<Cm����1��8p�~8�8�8d	�yE���`AـP*��qP|�9�sf�W��m�R�*�h9kx���:�$�/d����D�����F- �BQ�� Z��v����o��6���b,p����ԌL�.����Y.kh8�9�AFil�?�PWyʮ��0��;��8������/b����xQ��+R����#5���+��я��]��`��O?����<����j�k}r�1Ոܞ��`��͋�z1�p5��d��W�M]�V6�'� ���;�k��ԉ;��V���qQ9lT�鄯`5��sL�+ڶl�Y�N�����^���ƫY۶�A�r�t<��*�	.+�;���.I<�US��E�os>�V]���>"��rŔ���&N��%ɶ��7�"�rE����'�Źy�ހWj��n9��y�������/e����3�h4\W���s�s�t���ϵ/�]�奞��p:�ޒ�d�S�b���+ŊN�#7\�,��%mNcԴ+���{�e�d*��[noO^C��R�=3;ۗ��:��|����U�b%���BY�&�9���<��r�3��(�E'�+h���z��@a� 5�O#�D�|�wT�8`�q�~�\⇡,�ّ��d_�Ĥ���r�{�a��-'ly��6�f�,8}* �؟ l��֛	�T�U;��oR��1�e��T'�d׮]&��2<(�H����r^>T!5$��O����P0��@�\�ܐ�����ͣ;�X����d�/=�/�?��m���P\�@����%M�
�-����V��1�e^����;Q�����b���ȵ��;����~��㿝�W}�XU7{"z���0�\i\�6`p�n5�!7�v��6M�g���o��`�4��(x�>t�4I8���,V[��i�`�h�g�e��cHخ~�ym��7u+�rT<�m��F���T����ƱX�d����m�����2�*LpO��iUAX�CKӲ)�K%����@@�.��ʍ{���g��C�{Zs-�W]b=��-��>0:������o�����})�a����hS��K�t:�L�:�fSC��ܶ�Rf�Rzisz9ݙ^Z��R�x&_���k�"LriFu������{v�b���?�l�i�@�::��W�����p:��manq�B:=���K�Z�Z����z�X(����ҠJ;�� �ƃ�<�T*\Ϫ���<%�(�����*�9#��ܗ��Q]�h[�f�㷂��\C��W�[ao5�H��-��*���dP�#��jҫC�LG���*��B�#X�u������gooO�֭[5_�P�I8�q�$��RF=� r���)C1�go�˅<���9���������������E���9B���ч���ܬr'��,�V o�"[�ٻ��ۤ��;X�|�f�Y6�-z��wDe��󝛆�~��r5k ��m��`>;ۈ~�����'�q�7r���l�HLb�%����t�1`NM� `k@60 k������B����ș�fh4�&��e��4��H�����q�nj~�����\ G5
�q�G��ŬY�����b���J���y*� V���xྸ�J���l��<�C���\�.y
,.f^_7��'9�)����4 |�(��$B��<2�7(;���3��K�� �n����X�	�?���Ůt�����z ���d���J����w���'��s���x6�Of����T�oan~Kz9s���s�BW.Wl/
aZ�`2<�[ܽg�����6|���󱑑��kn��;{v*�ϧ�r�JG6����]�r��\�g��m��Tw.��Vk�j����@�ֿ#�ӸjuOXk���֟�F�cf,�0��((F.bO2f�Jc[7�즿<j��=_�Ҏ=j���\�o*���Fib�1�q�zt�۲�qZ�X2�Zw;�p]���2G�J$R0��h�K���5!P^����e��]�Qg^��erjQ�^���#�FellZ;�i���V�� 5>�f�[`� ���*�V�c��K^�V�����`^�r)+ɶ��u|j�殟r�\�}y?k
��t��o���?z��_(��̣���L ��NU���}�!�X���$��m��af#��P���;�r�˚`G@o�_3����X@+���d�;�m'��Ԓ9ff�rCyA�v����:�s�c��='��װ�6�ӕ��C������(���95s���`�D!W*�[��y}��
��$�>�9�Q�n���/w�*�zM�/P3�^4`�\/�r%/U�\�B�d�l�;�P�`�C���3;��W]���������S��a�\�}za����-�s�ҩԞL�0T.�Bn����z�}�l��厎��m�0q=C>y��Fӑt:ݖɤ{���P6SܒI�w��3r�|g�PNV*�x�TQ����ʬۥ$9c���b��/�7�c��a�S���9��JܾR�:l�	5Qω��z����n��'8�[�`Tq�qw7�馬h�%��lz M�р6�c��i����ke��B�߶mۤ��G��g$QWHB�vYZ\�2��B�|*ȍ�v��o٧�d��k�~�-�3i�t�tv�KOo�\�<+�)A���#��)Es���������9��q+`S���#���m�K�Z�X/�bFb���v|������6W�zֲ���=�[?3��y�{���O����B��s4Hphѹ�a��E߬��5Ȧ���6Ђ�-@$�]bN��)���`�@�9�qnF[) (�2'`q�����=�٨Um�kU��p�]�6��I�E"�A�%�g��V�秇�������ι��n�eݪ��y��\�nw�Թ��|&�`�f�R,��T̋�R��`HڼA�58$G���zT�n��[�����!>���G����A�z�R�6��nH���|�Z/y]S����}[��ټs��#����k~�Zߟ ���m˥娻R��C�Z ������5�� p��Tri)�V,����s���b:�������r��,�*�b�ꃵhm�n����)b��X�3�����<���EI٣IR�Qo��_��
C.�{ �p��x�}���jf�҄���;5����й�\rbД' m�`L�Kƨ1��׿=&7�ݬ�
F?�����jY�D%$��*�3Z���Eٽg���Ys\S\2;�,�/\���ٴ�G.^Zж��k��Q)���F�@X�	�&�ak�~�`�*�Z-��0�7��u�o󪔊9�Ƃ����Ц�޻�a�u)�k��������sc��U]�1-35�hi�w��Zj(]�+���(R��(R���E�#����Z�6�0�n+
6�*�SK%�~q�6
�`or>k��7�1�M����|�k��w����ǲ�f� 5p
��E�L�� �;Z��7]����c�O�9�`� 1lA��@�e�YqX�0�5�nU����wd�<�����%��I�պx�%A�Gbހ��U�DeX1�HH|h���J�Z�T�$%�k19<������1�h|��z������266���$��b[!�ߘ�g7..f�.����+՞B��,ˉJ�k4AX�. *�\^�҇�`���(�T`u�9ʲJ%䎠iHI�: g�!ĉ���P��]ьvĊ��Fy��*KQ9�Qrt�S9���ƣPo��z5���r�'�����o�1�C�j���CW��xH�4ދ��69t`�Kyu��y1^���}!�(������*˖�^y�]�R0*��6����\�8&�h\�m�+W�dvn^�e$'"�퓕����x@&�P ��l��ƒ�����M�ΪLn�[�۲�ʜq9r ⱐtv�No蹫�3p���kj��������}���/��R�{lA��+4��U�-8��]�$�	bF3t0}E0�ڭR�����C{&�`D��]�����m���jn '��nv�i��9V�OM���w\��A�����y�s�J��K-���=o|~z�<z2�EK��1Cܓ1s���$��I�X�2z;�sⓆ$A	�\r`�.ٿm�L�� �tV�.\�Z�$mѸxa���^�I,�E$H,��?"a_@�p��}R�{%�*ɒ�v&8��孇���ѣO�F]��x���?  �Z$���b�/��ݰ���r�-˙Lo>��̕��z��Z�x3���������gU�uA+e'A�Ш��?�y5x�LƸq1�N6�9� ,.�Mw*װ��.�?��u	xMKP���c�u�����j2:-�סQ[`��V�e|��!	G��֖���eyL&�%��r:+��%	��U������O�N�������s99w��R��ܽQ�^]4�)��\P���gƯ`�X̃&ᐞ��s\�֜��s4�\��>;<�]m�C�=o���?~��zM���K������ҕ�#orx̽�@`�9���Y�Ζ�7'��h�o
'ֶ�i�ڠ��6M;A���D��`�{�/�rZ�B�x-Q��9�]�n/�ck�m���	+&Fn?�����<^��6pL�����cl�6��e�
�j`�+{�셂&5�C�ܻGn��x�dX���?$�Wǔ�
����%%G�,�\^\�Djn������#W�h[B$ꗩJVf+�j�����޿���{z�mY�~�^ɱ~�7���K�`ї�4���L1�,�*C���m˹��Tjiczi��X*'��z�Uw�j��X�$2;T��n�O�����T�J����f���5C����ZoH�b.�LK���� �j��$�<�~`[��}��a�*��y`��O��}j4��4�e��=�K�>�e��]"���C�-u�!�'ڕ�o~nN�A����'r�]o�h�V�@��s�w�;�Y&&22>1-����&Q�>��%�+���Z��JUF�C���Y�i6��E�H�1�9��"�eg26�q����{����-��`�����~���|�����9�'�hX-s��iN���&ف�6X@v��Ws�t�u�.6�9� �0l�����l�������E���q�<Ma��Z.7�=V�uO�Ď�D��    IDAT�s���TM�$XW�}��X�X��l��N�p���5�l�Re?+��LY�k���ΚD0�)�,:I��{���}�o�y�Ӓ^\�K�.��Z$��>��-푤t�1.Sk�[�He)-��e�fK����DP�ޖ�z�#�FAr�C����;�n�������w��>�n��|9����l{.[�ͦ�����b>�5�/K��|>�U�T"�MRm?��)�9�Չ��{X���l�ZqBV9��ln����	zw�f�^G����]u	�LΎ2�:���p1�B�����# �P�X� s#�`j�	Ce��HUexÐ��v�������M�<M���}ޚ�5y���H��͕ ��tQ.\��<��Gev�(W�Nh+T���fQ�J�	��a�SƩ��l�E<���]�5>�-���O�ul0���GtW{4�q����vk���5󇎟9�������������[�9]ʹx9�V@`6��=ZeU6��`n[ݼV+@�\]�N�y�6F�����8�8��t[A���L�=��:1s�9>k�4��c�(��k`O:IZ��x�y�8�_qCY5�|g�c�A�r`_�:�s�<B'���`��P�m	@�������c��LOOa��h�^�+ A/�8�}���n�$VsK���|Zz�M��TjJJ����K�S���'ջg�gw�x�χ_�o�E�z%���/iযT*��l���-lL-gG���B6�-�/tK�b�nT�R�@SW�70ف�9F�jM�RBM��p��\0$7�E�o��6МV×��ұ��^�f��bz^�(��4��	:	pl|��gX������+��}��}p^$�����}�������_�*��\K�<��v�⤠��C[%����KcJ:#�a�s�LN�˸�M�Э`��V �Զ�&�t��V��6�؞R�X�9ٚ	��h��U��z~c��_\��ZS0����|����{f�R�3��cզ>M�����9�ae�-L:��u��4���5��� ۶zmE����`kҙ�t�1r^��l+��� 6W+�s�؟�[-x[���k�&��Z���m '�ӊ��oϛ��p��9�߶BCo�m���T��TF*岔�ޱ��NR� �$|
�{�쒻?u���dG�vER� 1M$^ͧ�"ɭ��*���i�.-�;_�H�%���
��^��<^����b@��)�7�e��=�{��vv�b�����>����ltq�ϖs�T�?W,v�ŮR��U���r���t*ӟ+���F�T�I���N^�V�G��Uď_whY)SI���Ţ�y�^����*M/�	٭,�S��3�ly��&�,A�
�+��m�-[�H{{����4�
p�E�$
��܂ԫ%%�A�W��f�4�e��U�xd9]�˗'������R,6���+���)��]���3�:Rӌzc����o�~,]v��3pm�e�b|^�o����ƣV��r^,'��u0f�;�2<���C�߽ޥ��`~��z�?|����o�׽JX�FU0Ýb�9�ʕ�vFnO�|�.�s�:��g���g�V��l��؉c���m�� e[�6Hr�1[1��o{p};	�Vr8V�����15�O����E�_��c��kQ)`l�U���<ًs5��51;�`�C��ZV�~�U����9rD<(w�}��K
�l�Ñ�L/z�<�ҨV$���Ź9)e��(U���H��-�N�JH{�#��&�UC>)�<�	��=�|l�-G�d�}��{�l�z����ߛh4��E	���|zq`zr������NMM�+We`9SP�nh�HSW+��$�b���˃zr�G��hz�=�lƴ!f�V-�nv�@���l��_e�
�/�&J�N��nu9��M�%���^��'`��!m�ݨ�%�H8X��n<(;w�ۤ��3�%�reJRi9xp���!�r�O�����ms�o8Z��QC�������Vo�6�x�mp���s�o��1���ɤ��3!6�����į�\�gT�)��s�����������9Z�!f�B}X� f�lth���( XD60�ͮ��$bgh���Z���nx�T˺Z��i����+�����e�qЭL�6]��xmK�?;\@ 5٠ƽժ����Z���`��᝷�K�Z8��A�sa+�i������%h�����:�LVJ�T�U)������G��;v���S�`Er��}���x|A����Dk�CA2����CDS��k� �BU<!�Iʠ/*цG�c�Ѡ��5Y�Vſy��M/���{��|o�h���F<�_u}^�4��3�C�S��x��ۦfӷ/,���fG�{�^1�Z�8��m��'(��`��u�;1�wX�P�S)��{T�˩wB����H=I��4\AI�-���+�3���u�88 }}}OĔ�=	���ק����C��U�o�/�����c��V��\�:�.y��`q��0��r�E��i6ַs��Z���ـm��,sp���I:�����ƞ�E7��B�u���)��_��/|��?��+� s�Eu���� ���i���bƥm�x��biA��4_L����� g��[�~�2��� �D
&��x|�~���m���-mj����Q�n���a[�t�sl6�75l���E�o3).L��r8狀�g��f�����WJ�0p�-��TC�>ؕ���DRM2��}����3��r����\S�)PT�n�X,"�O:b��B��e$S�K�^�B�t�r���/�%��H�x�G����K��W8 ��W��u��m���mz�M�mܘ\z�bw������@���?���[O�p�?�=��rN
��Z�Ŝ!��תʿ.P�jK��.���!c����f�~����G�9�5�w�5^���r6�p`@�{�w�w����l���iK&%W�I(��*��c�=��g{V���=eٿ�;�K굊���|�*�r��Uٻw�$�!9u��d3)������}G���#Ƴ�ߝ��y+��o�Z�o۠z1��u�#L9�� OUV;Mw�~x%f��-*����8����ɤ�dϚ���������=��B����I,�P0G�� ����Lp�خn��Tń/���*1s@Z]���Nz=��ϋ�֠��&H�nt]�X0�8�iv���m�s��`H�������-�a?7ǰ�@-*WX[����pl�Z��B\�=�Z$���xxorJc��z��E���Uf�FM���'��w�m��Z\ҹ�z���:yF_����-��6�˴G����੐ϗ�e�Ssӽ��tG�Xꘟ_�Υ��p�{
	�\�I�'([���$�+��eWU�UI�}v�m��dǑ��%��{�H�W��f����.��3'N���܂+�\����TK��N��1�
*�@�;g8��%^�[cȔ-؇��!���QQ1�0X���r7��5Ծ��΃�o[ww�=rD܍�,"c]���I��7�u��{J�ʕ��A���h������b~�n�Z��\To��tw'���f/�E��kP�Ab��a���
�i��r���Q�`��ea����I��za+?�|aa΀�`�#�7��%qM]��X30G\���o<�����P�8���2�����Y���jo31gRm���w�Μ���{5����&�_���mn��Iwj-q�x�	�Լ���s��Ǘ������-H	ض%O���,
n8.�޴���&���l�ߌ�����#��a[��{�K�vM��`��䲒/�4M[>�K��ۥ=�P��={Ԃ��r��ey�'�>5�hiMOge���/o|W��D"�����\�Ie3ɥ�b/]�|���������t�S���
��h�M����1E�S��x@<C�'v�~�O����������l��c�g��5_���_|�����|di1#��K�Վ�&]�r��9�̳2;7-h+��QН�B���%������v��<̱)߸���Kɫ�7�rX�ɶ����j�nv��h�h�Tj�1Ҽ����aؚDB ���H����[4{_�A"]ŀ�Ԥl���.9{nV�f�XF��O���D��̙0#[>k~�6��2���e�7v5����!�(�8r������#~��o~�Ʈ7&��K׳������O}���~���Y(6�n��[����
,��t�D���n[�EZ̴Z�{�`dO��Ծl�0� M��u�hF�$��X;�
����Z��[A�琮�V��jM���r8>{~譠��F5�
A��Y��7�5;�q^�De�r��v��p��K�S��c�F�u����;i�&�y}H����¼?��֛��J������][�td�֏��؞��?zk?�䩞��S#gϟ�����7_�ridyb�'�*�o�u�H )]�$���]��%�s���{�f�MG?�ig����\�Ǯ���c����}����kf~)�L������v��_x����N<#c�㲼��D9d����q+������nh�5���NBe����SF�l�d\\�L*��$�1��U77�u��ׇ�+��+X�i|
�[����6yӏ�B��|G�2���Y�����6ٱcH.^Z���Y�BJ��j��̑� W̨.yx-4�o�ؘ�����̶Ln}�<��<�w�RIǅ�<��h�#�/l�������Q�����5b��G���3�Z(5�o@�Z-s��kfb�	N��4e[���u��:��ɵ-oH[�̨��w��e�1�c�	�������U����ÎY��3�i5�X���o^��f���L�#��9?��ٯ�׷���1�ñ�:fN��ʷι=p���9x�K��ƴ���ZRb�޾n�����j6{[G��NN�L�ɓ'e||\5xW�"��n?~����x㝷~�;� �x����ξ����N����/+O,l�(y[�]�]���C^��n�6��<?pp�g^v���{x�s��}֏Y����<���w<���13�N�u����l�� ����'���r��)�x�LM�H���>�
f�2��z{p%K�d۔�mQnvݧN�@4�𜡯;b�9 �t.��dOP��M��l��9M�jфW����uS�z�^�HggX~썯�P�$NW�"�J]&'�djzV�!��۷]�'�dllJ�5T� [r�+��!�!�7��ZlE˞ 4X^�ЏmC�y�E��"���y���s��n��y8�����3Û��#8u=kh��|l,������ϝ��K�2� �3f�8��� ����t�r	�|g7�����t�ؖ2�m[�j�j����ok�v��o�1�W�G���fg��*���V��Ģ�� ��]h�Ѐ�$&�P��s�J��1����Em���h����!0i�~?vB-s��A@�X�9h\��T��>Ǳ==]�9��I��Kgg��a�����8� �_ٿ�?���7��ѣ���%��|��Kɓ'��������S��w�;�.�p%�J�Q�l�+S��L���#�w�7������O�\X��?�3�O?=z�m�<�����^l/��277/�e��=��'�y�+���Kru�,,e4�M���򅌒����+�7�l�GҨ�Q���7�)�!r٬�8�~���Sx��)�=5>����j|Tk������x\5�O��4�bu���R7{��d����5�ʆ�-y�g���^���4�9p`�����ҥ1)��iE�m���)������Ƚb&�&�9���[��B���AD��[q�F�mDQ.o��[��Gd���o������uɴ5��ә�}�G���٫?U�����ue��=Ni�7���%�X���񶀹�%�8L�m�����P�	`6���М�I;��� 0��n|�t�7�o&�K���g���(86Ƹ8MT��]�HL�� ���� -��+.2������n*,�}��P	�'�6[6Vƨ<����-�)ULM,4z�U�ؐ&�%i�6"��D,�C�}��׼�׏��~�b����y��ٷ-��������T���6�[�р,����Ҹ,�*������k�x���7<�R�~����<�����o�����J�+K�����ؤ��K��xXR�25=!�Y"��Zv�6��dx���#�-7��e�;\����P�E~u��S�Z����rQ=�bAH�\���.�W˦M,ø�Z�r�p�#�JZ���ؿ]�+�����/d|lF��|F�9$�\E.^�*���D����幌�_�\�$lI+(���6P.�F��F�5;XR6�����^z}S���z��j�\��W�ߵgW�����̯^�����}�/ϝ�|SӂQ}�A��9`;K��p+��$"�@Z2�5�����"x�Ķ�m���ͶR�2qi�{�.���q�8ft���(�e��G�X[�_"�a+��m��ul˷��c;���%��K�p�m��~��r���a���`k��\3P[��C��1�bq�x�c-�V�Ve�M�YQ>�*�7�N��K-#Ca��a�'n��ȯ9��%�9���S/t.��r��S�q�'owM�<h�
��j2"S�\�/�`&w��n����������ɵ���Z���2�x��-<���]��T�x%jh�	0��/7�t�ҡ��sv~^|��Z�P�������2�� ��0B�V�<�d:�gB���\�tEz:;dhd�\�pNr��&�A�`��x������#���=�� �9oL�V�6�˧$蒗�rT�m����tNΝ3���LJn��F=���	YN�.�&�`Te��\�bI��0�!���h�tx �Ú�ů�@�`�(�F��jH��nT�]<Rq7�5jnw�0v{�5��Us�=u��Ss���h���q��n�� W��v<nɺܞ\��(��]�z�%�/�s5jiW�~����d�+�ka�,��6���?��+c��!h��~��^�=~'va���q5��H��y�%F��XeM�r��>ۅ���x\Hta�xƽ�}]P4�4M!ȡm6�}�+���1Ӓ�ozx}�M:�c��bia+xW�׌�Vjt�:mVm+��k���/O� 3XyO�������g�L*d�:�E�\�B�����@����Bl�ɑF���zM���9��!�n���[o��W��7~����x�q<򩯼��מ���	q�����L��Sr������ҡ���-o}�_���v�������3����ɳ�����G?�¹�=�_���/+P��/;*]I�����V@3�rU�1[ML�朄��vdCXKI�r9'���6����?(�JI���3�.��R,$����؟0з��E��;::�c���q$��{����/LK���)5�喛e��a�\�P,.�tA�}�y)�RH-����d۶�r��΀�	{��[`����s���5�[�E�R�V�H�j��;�r���n�5��6�K��;_��Rnid�>wE�W���e��S��ՠ��{��Z��!�P��k�F@�,h��u��
ի�Z�V�$����-�jk�[30?wnf�߼��L��P$(�XX� �K����{ʊ�����`c���u{-��uL�ֶvmw46�m���gA�.cn0�-���J6.)S�a2�#��֬��G�"���8�	)|>�펇�i��{q��y.=Tn`
�����Ί�j�B����U���9/L�a�\]��=��͐@ä9 9��A�z�Ў{oy�M�|���k�i�������̗�"u���.wDKx��̺�r|aR�Ѱ�m�t嶗��?n�����o�2ŷ�?�3�O0/�0��K<��s��������%���c稌lT�d	��9���WOW.��}�����M�LV�[�?.�d�9)��0�\S�C��}�4N�;��8�{�+8~ppP��>���W�y�e�+d�T>|����OK�ڐ|�"�3���V���妣��4mvfJA'�"�P1�W�sԼ�����]5I&��D$xO,�X :�����<<�V�V���~?�Ś��S'.m�������l�0��င�a	@(
�͸D}�]V�=�mZ}&q��B���k[�6��������+    IDATq��(�u����N�=�l�� ׶��LyZ�|�&�3��cl��8��:��`K���^cG����p㭀�U����7��3\���;&�{AF)������\�.�Uε`��]-sW]��zﭯ~ٚ���Cgb���_��_��eo��j0(�y|�\�g$��.#[�|��w��{o{�+���a��>�3 C��|����_��R�����t�d�{Qz��[�ett��ے��ވ\�%Vk&c�␬�Ngd9��t*�r!�V0/�*�i bX�HF��޸��a�Syg���Q&&�W�͛7k،�l>��\[���z�̵wt�;`8���9	�R�#񮨙�)KG,$��v�d3K�ͤ�m��-`A���x�A��Lw�ԕ�ٕ��כ�Ձ��].��'� ���?��Ž��=�����d�/;��H$���O��7@А��u�W��M)�;6��b'��V��B���~2�[��d���&no�뭖?���q-u�x<zA�?�2̰���F�}��=�/���Fk��m�&c�,��+�%�r̨�l�|G���1���V�V+��\�7CxVd��0>u�
+-P5�fY��N&[�J�.:��kr`�ֻ_��[~����k������v�}�*]�;py��	�����yyzrL$���.ٻk뽯��;~����=���_���|�3��Ï=�g.�Z��4�$0F�J������l޼I�z{�]�}TFU@�tW[\LI!�x{FSU�������`j�l�tJ[c�n޼�3W�C��>R�"���ɦMh2WT/A&�tɷw�iS�H4.�bQ�'g�K(��T��f%�m���|��<O--H|�r�c`n�8��FE���'��P�Oww�}�s����5�~�����/�w�cmQ	|�f�6L�x����(���%c1�ڰ��s�en�9A�mK���RlEa5�;���~�@�w���Ǳ�������xf\.*��m��`N��mկ$�UMb~�lu��p(U�S�{���eu�Q頇���J*?��r3S#���o��`������ߣe.��e�k#f��Ua��+G�|ϫ^y���ڵaq-7���O�?��O���GO�L�7D�F$*�!�<z�d�n	u&��+�x�m7��[���?��������˗��y��>���\�eP�/��R�P�J��Np+����V4h���ݭ�bŋ{�PR�-hqR�����/���3g���dϬ~V��m�ps��f2(7U�G�*�!C�ی�u�{g�>��`�c�h�S��:I��Y��T���b���=���9&��{�]���yQWQ�Uh`g�:ʣn�Q��qw�T��j}��%���B��^�0f]�5���҈Q���_:����-n�g�'��vJ�7��U��9+
������<���՘;�n����n�5�˥V��ػ�^���7{�E �j��7m�V�9Ҫ�L�� G:U�����UpX�IX�95	:*��
�ԗ *�asrU���k�[���cΊ$�OyO>l�}��ǣC�u�ă�nc&75I��au�Vه/�l۲�<&R��r��˙�K��<���{B�r~�������B)�9v��?##_=,��&7�.�^��{�/:BFL�^�J�\ޖ"=��9N?����<̫<�5�v�iĄ��28�f�T���Q+?�<9295Ք����t«3Z�ܾ�e��p��6�.�6ǧ�/`���j_��%�������b�d�:���T����q���G���CΔ�I
��	Q��i*$��.��5��P�$'Q��Y-���8�ԇ�F2����������*D�vl�ՙ�!��׌.�V.������O9�y3%��p��V�b��ɸ݈��{	��s|���:�
~��#v�<K�Q��fJ�&�b�㮝�>E	�Վc-ӓ��z�7OKMF,�5��+@��U"JZ5����h����Q�r6iKt
՛!	�h�\o�t�r�Kn��6^{����8/	,�o>Y�|������@4'����@'zE��7%@��# /���W��V~��L�>jW��6�R;�2�da�1�Ǭ����n���է����F����X�����x�9j�v��r�R��!j�~�'���ۅh�{�#�<*y��U(y}?���r(��/�N�w8���ϫ&wF�*%)��֢؜��OAO�S�c�5���ŋ��8���}�X�n.�{L��6�z# 5�(�MWk���+��#^�vvQNZ�丒� gg�a��Du�6�����On��K�����L��	��N��K�,sJh���M�4��YzC�6\�׾�{���g2��U	���G����+����@�*ں[�`�!�"��\;h�Eb*#��s���4P�������.��� �]��x��_���z���1 �Ih�:>�R�a��xa�J*\�k���Ž��ޠ��'[��df��9�w4���k�cj��(~dIM�����Oj+	���z��d{Cp�{���<�p�e+�z�ǣ����Fj���Z'��<�����ن�_���Q]��н��|�;.(FI
�vN3hf%0��В�/�fx��u���r�wv�TRވk�6a�}Ɛ��8W'�|�I �Lj�m~َoc�	ku��UN���Ka6�ȸ�i����6U��]�B�
�(��e���LI��q8�e���P7��Y�r\��1_�M�[ 0��XїdͶc"������sAZT+m�b�BT�c|D��]M�7�Lڵ�����߅����1J���{����F!h*�����$fp#�w�/��RR��!;Ѷ�5�!����=�E�q�B�,X{ޯ�(>Bu4�;:�hO��3ь����1>�5�@��8�8�����i��?kM�K�v�p��4��".
�(�bM�̰I��D�[/Q����{�w�"յ����a�����_[��~w�������6�>�C�0���G3�2wu2�B�	���:Mڷ���h�A��vF`mI��G�L�s��r�?ik�8��Pw7�Ϫ]2,�r���7�-/Q%�>�,��Oy���/|�)~��I�EO?��ǿ��-͝#�ޘ�.
�S6�	P�~(�I	7o?rq��V䮾�׵��-\Z��7���ِI�>�Ӵ�׫4W
ῦ�K�(��0��vѲKp8l'd2e9�:e�ޓ��r���.�RDD��8���6t��ȡ�[H6R��h(�+a��K���ϭ~[C3.�t�ۯ�J��&��D�6c�	���i��J��(GV1�y��xd]U����k/�Z��N��1w��[�����8s�H&_��\���vu�x�c��V��&"a1s�M���^l�7�h���Ќ42=��.m\��lf��B���۰��H$�KY͗/�X_AI��0k)���_4���X?D������P����\�hgV�Db�za�I������L`k�"��p� ~���\,^ϡn�a��^e�����z���:d{V�g�v�ٻ�<eY�2S ���)2 �e"�N��(4p-R���7:B�w�>���� �J�&Y�W�麵g�ޭ��!��v5o��2�(�x:B�L<N���`;|n?<�V���5<�=��W��"{�jIw�����ߖ�m\(Jf@7�j%�{�QQ��}`nEX��+����-�p+�E��0|g:u�M[��{�<Z�H�)�$��l�Q'���(��NERZ�Z�m�xLWF⏶R��$��x��|f}ėsP��|"�����I����;s���17�:)����$�Y �<����i�N��.�������!�dcMK:ԶV/w��?|s#qH�b�������Bj�����R�j��:�������7#��HOxx�b
�٦�q���޼x��=⡹�ٖZyJ�G+�ԧ*��V�M[oο�Ɉ����4i�*974J�D�ޑ/l�/���:�N���Q���������ˇL���ʧ�l��5.���؃7m������B=���L��$���ѧ���g�w������G��Ϻ?ϟ��zl?L�L_&���&�9^�c9���\���i>�ņ\5<�á����0���n;����Ӣ�:JR_X�)��۠��V{!��ð�m�g���S����#�o���`�;z���H��&�[�o�@�[Z���dg,{�T"���3���bH_��,��$Qvo��(���
����ze�!�(�7X���[O@+�~/���gm����w�������[��t�M�2E�ŀ�B��ũg�9�����N蟋	B.n��ޙs��)z[����7�о�,?�! x��g��;��&QGGJI_p~���t�	l
g7n�B:]3�S��X �G*.im�v����aq?5.{	�n�LJ&a:�Ao�P*V�߽���+�����o��'����	Պ[�߱�S.���d��2�j<�p0��ҟ�-��L���Ү����8i�cj���I��zr_K��ع*�5���q9����)�j���3�Qww{��iJ~?L��,5)�8��]�A�L6�p�[�6������9��|M�v��}��Y{#y�������O��nŰhv��;3�����!�z$
�5uc�|��}8F���
"�������m%�5e�pf�y�%`�h���5+���H�k�}�b�{B�S�Y�X��i1�>t�i�m�(��e�4U���r�2-�Z(��W��>�\���0cc�����U��iGf姈�k�t�(�����[����
/D����&z���B{z�#���55�}/�{=�Z��"��`.�tU,��|D�S���ͅ
ǢrD8���5�Z�� Z���D���ܱ���:<MA���im��]�M�B __�ŗ������a��,����ع :.�Ǽu\��h>k��voV�j�O�kiq:���7Nm�âl�7�������a���8��Q7�d$�i��j%��Ǝ����wh �^~-�\4�6DP���;��1���s��Y���������o�b����OI!�Ͻ��ާm��+��͖5/�B�N��Ǐ�n�Nc�ɗ㕍Gd]����Yg���+��W�ݠ�#b��ۑ%�>&X��(r�O�W�2��ǿ�7	e��y�9�TÉߏ�a;`�]������
�!KEEŌ!<�������\v�Z�5[��Zǐo��b�Y'�����X�׾�O��»^���		�\�Duks��I�e�����S�۷��#��b篜�_��n���Y�I^?my��z\),�:*@��������q����.d$���]og/�O	���	��e\'&:���<��)d���^�)�T	�&d�k�va��-�	n0�௝v�6���`�I�g�}?
u"��g��j��"n�(����Pky�j��8<Y�����-�C�}j�?ja�7Uf=��cw�	�j������
 }��=?��ei����L��	��j�B�P��-�x���Wk0�R"�W�CN�G+���F\�`ܦ�Bl���t~�h���)yx�;��7)1��&vxXo��;��%)���F��
'`@;����{17Q���o�ϫ�������Ĕ4�2��ƺ��?���n�WO�����F�B��v�B	_oU!cR���M#y�����b�?IK3ǫ�Z������!<�G�|k}��2m�qў��H�4��m��;5���L:��o����W��	��D|D�>b +�3�\o;nWi�]��0<==��*�������Y�D���d�h�bE� �뚶��ĕ��.֋��烏4����ō����S]ɷY���d���Y��F������P��c_�bK�@�K��zzWI��z~ijy���g¡8%|P��r�hi��w&���7B�����rE)L���a���f�Ө=}���r��7#���y�mؓ%6Ѫ���^::��o�-.��d9ƿMH�'��Mjm�+E��-��T�ЅĄ%J�шd����W?m҆�tq�'ʹ��؉�6���S�C���[�J!�ݨv	ʀ=t.��}�n�1�͏M�Nh��!�
0�#���NT�!_��Be0a2V�8���r%��Q0�\��P�]VN|��%�|��*����=﯏�.}�z͇�Ț���9��{1���T/�'�g&��O���$�`f��V����c�N>��o�� �H�ce�L�g 	��b�l�Qj�#���F��G;Ix��Q+�_�o��e��2��a6��J��4Ͽ��99��8J�H�dE��Gl�%�U@�e��%�#k6�B/�A���R{5;''�ʎ�"�r��Uh���<���
{���؆{H��������\�������VȂY�Q��F��\�4�&h#@��O�E� ҆����z�q��ƑQߪGR{͕C�Frz7�PȽ�E��3������Ƣ�r Ô�D�@��"�!����*�q�)KX��u55V�mP���8OO�8�W�s�!t7��H�!r^�������a�j��LP����{��m��hkm�8�!y���I��ɈI�2@�,I���� '�#�d �AҪ����͡�ζ��'�5IZ:g���m��cɞa�&X@D�+�wp��^��Y5���DCh�+(�~y�%^O_n�P���	U�Օ#_s\W"`���������nd�Zja}_�Jx)���GV��5'�deT�K�z��
*
@�������Z'�zx�1�f5	ݱ�<��XCN����q����$�#Q��r�@�=�M*�����J�Q�����f��,��i�����Ou�3�E͆�{"RJ~9�0s�u�o��.��4�T��^�j�};��'+:	��ů&��-��nQ��z��*�19E9Y�w�l<����xT���r�u��?��-V����E���*��{E���Z���F�y��/G'z���r�Y��3����Jk8�O4�r����}�.��h䉢�G0�+*�}r4"�@�ۤoX���@ПXTik`@��i�������@б~A����@��B ���ܵ�a`�s�X-R�F�s������
�WGD��5��I��S�a����
���@��t�0� :����^T�F5�[V�2H�RR��E�]�A���Y���&�"F4��R�lL;?�+nN�٢�A��2\څH�Dق���m��[���g^�-���r�,ĩS�ֹb"æ��	w��)Hf�Ȋ����ֹŅ.���R��\�J�!&����F����"�����F��.>Pwrb�3���IF`3�Z^��Lf:����|�4�w̧FxKM�]�Rw��65"�!�����W�	�/t���,��?c���H��Y�J�wӴ��
�X�=��}d�����T�ut#�E�*$�.~CG�(�8�?��]ah���W{�LO7�'����\#wH{����t�@m17lX�������+A�W<s�6%H�W�@;'��Z�X���m��"%��~�v�;fy�[,��x�z_�� ׁ����״�+9/���f Av�}�Zt����ǋLf\�޾jg��5���_�k��0#�H�22%%7k��c��04��E����j�D��ݱ�9O[�"9��-�>j����Tpna"^Wz�C�i���f�xb��&;��O����)��oP���Π���6�y� �2��8԰/����	�ﲊ��֢�G�pca.ƾ�B�wm��m`A���{>(�֑J��;;�8��<�� �����P��0���0�"u�5x�!��������ff�"�e���+e7��^��0����g�cac�w(}�Y�f��δYc�*}�-����cje�q|���*t�S�$ePΛ>�+%%�v�nw#F��X�m)���[��ZA��\k���K���3��Ý}��A��o��/���.0���O�I���9Y�2I�f���k�JM�#�֛��)�vuZc~�����F��������JtR�7��Hw�k%#}���]��"yZn5�f�Q�vN<a�M�,�Hܹ�ȯ��6��,����!4H.��a�k��v�c��j�o��3��F��H'ƈ��یެ��T�&�eݷ7�)x2e�I��ưQ�e�^�h��t����H�0 q��V���؇?���_��^Ќ�M��]�wr��b�6}=j����ﱠ��	>���3�9�*��u�����gĖ�\��0�Ɇq=�(-��;v^}b�bPŐ�Y_N����<��Ch� �Vzn3V��/�~����MŬ�i��PgE��hK����8�#$��祛�jl���á�/G%��elS  �H#���V�LGGG<F�V��{�Mb�(^?�� 	0 4�a��*f�2���?UfF%d��R��a����d��GR��_:'�lv��'s�^���Q�s�>�Z]����B9�,����Z� .�4��	��\� �b���;����_}� :e��n�=�����>[������bG՞5�9�<�o�\�+�u��ڊ�KGe��D�b���hc����n��TJ�.���J^�ܲD$�S69�r�Tu[CJ@�8�ӢwYJ��Y��#4�GF@���2�zGd�F���7�Nt�銘>
,�)HS⦤���o��p�x�u?f��c���0�e�env�խ���N�6r5H ��3֝-��`.@^�;�^	�y(��o�*�v�S�lmw��T�/],�/?M�nz���Vt�K3 Sâ_���m�?��UQIf�:C�G�e��,��<��D�z�xk��X���n��p��*ԭ�ú�=ҙn������yLb`0]Yo�w�{o�<��m�+��8�`-ȁ�j��s�DY%,OfW$�� {�J�O\�`���&�8��\��f`��3��Mj_���=j:ō�16�Ӗ��Ց��T��w�43]�iԓ���>M?��뚌'��y��8�
�J\:^LD҉�2��8� ֛�QA��(t�G4�X�<>�_�'?�0�� !���=��D����(�c	��<'����r k_Sg�=�c�<�)s�f`t,~�	ށR(�v�X$b�2Bu�e�c�әL���o&j��PA �o�h���b0�o_kL�/��-���T%k4Ce�sg�Y��gC%������b��7?��>U�u�(���`�J��T��7s����(&1Kp�<�f규�B�=�?�*3��o.���\l��K�����C�j�4o��u�o2��W��ra�Web(��~�VR���D#�t"_�_U�{U&k�:���D*d�/��x ���M*�n�軍��>h	������Fn��b�z�.��ME�t�ݖ ���ܖ�"��U�+6u�L_]��&ߋmy:	��m�'gO���1_m_m�c�F������VIa�%� x�1���
`�.���i��H1��rﬄ��� 7��@a�b��  <�ܑE��̥5��g���a�ϝ[{�෕	Ak�,��c<a҉�\�+�T 
 +$�"����*�m-��#r8�1 n���#>�>�E��VP/�Y�QǙDy.��<����GZ�����e�LIq�3�hV ���l�2E&7���R�bʽ6�����+�+���.2��B()}�NJD9B�����M��F95}
��:ĝ�^��C_0�<&b-�t7��H�Iٯ8	�4ż~�r������{ixsʪ�:��|����Q�'���F��<X;x�'yF��9Cا�>�f��ͦ��9����/m�2Ӵ�b�ڷMm	�e����櫘��gn٢x���Aŷ#1����M;!'�IA�?�H�3knp6�o��׏�_� A��^ ���uV�L3�Tà~3#���;�)K��Q����$�D�L�fl���LrNC�9.��<6
P�L�X���	�*�����;{�7�5Ԣj�tv�tu;�QG rR/�O�����ڰ^�h���N�^6�f�p.|m�J�Y�u�O�sy]�f M���Ac�J�Z�
l/�2.���$�{u@޲B!T�!v�*!�l�����P�!ym�o���ʪU�GX��?'n� t؄��|YiG�'X��+���C{I��oo��-��зM��(�CKx����ˁ�I/�pe^7����^$�V���!I�����2[�K��������?�OJ��$(��myy�$�"&/}��J�#�/���4��ڿ=�n�[J�UP0�jLV0���5p1R_p�eS�5tސ.�4�6_m����`��U��K��k*��lp�+`eT��
���t}��ޠ����4�$�o������]Q���+��n����9�i�ד�@�ɉdy��8~��*��f��`�݊��h���pw�|��dA���^��VO!i�=�XDӹIC͒��
��7L�х��NKg\���)�C�n]��{���'��V��JQN%j͔���Z?�p =]�����N~w���j^���g��t��@q���T|�0�:������ۢ%�C��G��F%'�j�	����C���`����RF�N�k�G�x'�����E7� �Rǉ �~�ESQ�xh��AEm�D�o��몼��c�d�C�c��������I�Q�xܙ�F���(ރ�}��L�1��ę�du�ӍmL/��a"��t׎<*�&��_���Y��F��
��Y�op�}Uk"ڈ�t"�rc���6^��g�mz��ʀ���J��0n�~ꅭ������FkN���V-�"��z�'���������P^������Bv2�[B���6��:�'�,?����E�K����@;z�'��bc3��#�`Z
C���~��ǃߪmp{�\����,��FiUNYr��m��7N�|z�����6��E�j*6 ���U4��}�/꾄�$�j�}�{z��%��9W8�Ey{5h���>���~�H�[���#  b��=��U kC	��� 'Ʀ���*ؗ�����5ۈ�ڍ�}�����Ƹ562����mWo�:�Mw��Y�<@e4U�)��z�ƺ���B_�+A��=�'6 3�'.�����Dxك-.�A�&N�1��v��w�I<!F [ƫｿ>kB{�.�I88�6��}���8�l�wM�o璁���ߺA� >�ƪ����¥�6JaKMǕ�����Wm=�A����������i�`�^��Ȏk�M�w��22Η�%�矡��y�DN����b��0|����4�wo/�:Q�x�Ԗ��z�� Y=D@�|]�.�x����Ct&~o��n�X[�ɘ�&ͻ�s�s73���ɳ%ߊ��QL���R����_��h�:�|-�׬�!��m��nj����6%t+�L�ސ����;GR��� ��e��/�(��o�.����j�dxqB����~d~����0x�4k�g¿�y�����,y��������e�"�	�h��i`w{U�I�4��P�S�� ^KG�v�,��({��G��)�4Aދ^$hė#B��\Y!<n��o}��©�����V�9�p+<k*�V �7�G^��Du��J�W�vƤ.g�X��k�fiE���J�M�vm�2��a����P�Ƣ�[�)��}���Rc	����0�f�䘈�2 �#�E�������/�d�	���G�G/Dz<�U�m�"����Z|�X�@��-Ȉ�"���d��=�#Da����!��x.�$z��o�r��BaP@�G)��:���	�;\o.t�a�W���¹5�D0"��5�_Z;�f����l����f�{��(����i�I�㳩��+g���^� �P�dh�)L����j��l��x�JG�>�n�Z%��j��X�r�F'y-0�,����x�!ɿ�e(u$�!�c�󊈼]���`�m��>N|1KQ�v!��l��GlT��c��b��y�?�Fش�trB������u�����]���Sȗ�N�[�����4��ڟ�h4� ��?��}X���]�-<�0Q7��(��	�s�a��[6ц��a�����@M�y$�v���, &��*Q�U�:�dԭ���,ۗ�� �v�#e�]��^�H�����o*��pz�=9����QjP��|_`=�"��p���>�|*��W"n5��c��#�G\��M����x0�p��-����V��k�@4a��ཨ�3�ʤ[���X��x�~��K�Nqe����� 3�L�uF��JZ�}�E�HB�������Y+Np�.�n�����=�B�_1�����AM*ljq��?ĂOP��D�Y^.PJ���Iz�齾�1�m5��0{zlV�Ns���$�f0�9�Z`*�K�
o�A �m\Ӏ��
�?f����E��(�	���~\�I77��W>t�gU=�l�'����U
>�Bd��]}�L�}�ֺ{oF�9=V�~z�Vz2i�l��N|�3b �K�(�s�-&0�B���ޠ��%��軠	�\9'@(�y�6�/���D��f3TN�6Cӳi�M�#C��Ώ��I<dt,֖e�A��7�#Q��c"b��i�n�m`C�����>��m�!p�w !S����9M�y���������
,�3N�ζ���5�9��Qw1��p銨j�VN�E8h�g��RZF۹�ԗ�E���������]g�}���xg{%g!7Ó�|3'��c��z�n�7r��M���9��D�}&�<��0��G&��ʤ�{la�O,�DbX��1�u:L�D,�Ԙ�X�D�w՛����M�>j���%�=E]ږ(�l|���G��S4;�etg�X�T������w&.�T��@�7M����B�pv���©�9����vݼ�����3)`	���cɎ���Q{�?.=6�ME�*E#�6�'����7'~���3
ov^���s�/�N�eL�I�1*x���P�?��%��y=��"9�9�~�G�
d�ڊ���Q~HbA��f�KM��M$��z� ��w�h3(uؙ_Y��)N�� g������mӊ�ԧ�o��T�H(~�b�~���M}�˙����,�~����Ӳ\X�T4��/�y�c��צE�����h{���5��DSA	��=�jce�Dol~��Q�(z�6P)�"��5�Ya5���mfa��g �����2�nBG�Z�G�|����78r�"�HH�ACX�L\1io��e��F�J����gf4>]vtt<���;��"�Vg�J��]�Pۨ�7{�S1�tzB��k9[[�`�S�)�]�Pc�$f������|(>ܪ[�8+�zX�/��� ~�ێ�y=�F�9�#,����vpL�/��~�wJ��,r��O3O
o��+ ���)��;��^^�!��S@�4!�\L�ؒTB�qx�HF.Ҷ���X��1`'m:�����c�����&��@�������G�u�Lw(��h �����$���]\�i�^��7�����ͦ^e��+�ʩ%�?$��c�3��;�P'�(���ӎ�3��:���Rズ�_Q4+���7���m��J��BM0/�go��E� C,9n2�x��X0��֞v���T�	��xk�,�����v��r*�q%Iq�@�����c�wؿ���G��~�ݤ���}�B��Q"Y�y%O�Y��:������Us�"�g}�+��ܯ�W���A2c�%���Q�s�OϪ�jK����ڈ���{[���6���̂�aWW��*Y����+mB��5��� VYz��#y�5���_m�W |����o���4�)����pJW �����V2P
�}�8�AT�M�R4�iG쉨-�����o�
�Mjj\`g�e��>�U��(�}��5���[��!���	��F'��__h�J�������a�7��X��9,��c��&�DD��ս���Db��$_�JS߫j�MlK5�bT�n�����P��;t~b�r�&��H\ݬ�t^�Kv~i�w�O��*��b�S���^�� 		X�\18�f�:�wǦ��h�Sf*�ok'	�Tc�r��*����B�ꁠ���	��C�H�O��L�䷶M��-@你ʡ�`�cA �3���4$�g��k�G��<̲�(`�����B��J&۱	�A��.(k�l��W�����"���������^�8�?u�����i�w�v��/�A']( ���կ�j� �O�DD��H�v����^��j�Ȱj�
ڳ���7�hF� �ɴ��ë��pzTx��!�.!�|�Zϳ23o�!ϵk���$�TOb�P��GE��#�?�4_�9y�'v֎`�vs�L%a�"�d��}�2��eG����A)*������0_�j��4�N��W��k�@�)��D�r�}B�	�(δ?x��߈X�$Q��X���|ÙGe��q�Prp���-��2 �D��B�6��H�[�_mv�y�������qɀP|���] ���H��	�7י��&��x���ZN{mC3f�y$Z��q�jk���p `J@?� ���]�
�V�0��Ac�NZ}lq�r�G����3k3�d�'}_ޮ��<�g��1Dt�Vp^�O��d�_��*[�[<��:'z��=�g��O�&z�V�so'���T�.L�d�;�c���X*����ѩ\Fȷ$��
�֝�L�Q0�4*9�;�&O�7n2J ����D����t�~�Ų���H��� Q�Fz5��� PhT�D}�㸕���q6����ҭO���vY��L�w��h��s�=��r�z�@�_>���r�ti;jd���J�J����\G!ɖ�L��@�o6]A<�ը�ٚ��wi�a�,���A��)$4ϼO/a�g��{k*l�Ti,y�.e��bT/Y`5I%f�dmUBAb ˋ6ڷ�9}7zn
�aY�����$`��ܿ��"� �L�(9\&"��¥,�%�����Ce��i�k��]�y�T�߹�*b���ޚ�(Hiř�O�?d��� ���:�*��Z�|��5i��ä�W��t�� |��C�ґ�5x ���� ߀���rnhkw���8�8���
m���+�p�_���E~yfD�}9��2k.��h�(��-��P.���ʠ#
�&�`B�������p��?�Y�#N��2*��A6c�gR	�������6�
Nw�W%彰�{7�p]�ޕ�/�&�ɪv.���
S�#�&L����~���[��q1'��\U�jO'�R�J� ش�A�r瀼z;�1_����^ ��_P<�	Z��t��Ñ$J��0y�<0/�.Sd��0�`���Z�}���3�a~C����	����75�X���P�������̴W�?��W��|�^��"�Yo�ZE�gb3jI��8tڈ�sxF�P�1���A"�8D?��v�s��z�Q�t"���?�阒kG�ެ�����=���J�����\1�6����@��?�u�;����F��PȜk���D����>�ӿ��/��T���t^j�OP
(]E�W�7�?;isN�c��=@��j��39���QM =��.���P�n����&���ǁbK���oS�i��7���&�l�WoQX� �G���w�P.��WT?�x<+�{��)�\���]ZX�
�3��9O/p1L��T���B�b/B\��:�4��}:����f>ұT�Uzb3�l"��e�<�	��Vc�;�2�NY?�]���F1��I5�*z�}p�H+WG��5X(6���y�x^��'�%6O�n���I�\ƨ	�g��:.g/iL�O�swU!���$��	��kA�ߊ�˷-	�6���z���\r��M�m��9�f�d�����;�[��,$s���5�0~��n�*m���nޚ�z,�'P�p�^�7?��m>ĝ�h)6�Q�3L'=��S�o�2��X�XsB[���Z}(��Z*B���?z�g��������1<<=���]a���Ӣvw�X*Ydr3s���+����D�q`Z5��
<�|u
����y)OKk���`'E�P�_c���:�n�*U����v2��tG7\|抯F#��h2Y�����U!�\^ u��zѦa��t���ONT%��m��/'D,�i�!)�ʚ?'��Mu��W�q��}���Pzi[�!���-Vcmx��f�j|��'g�:���&&^6H� z���`��H��:E3�|T~�-��th����(ug��H�~���^z��B>��}9�!������cd5$:���7茁�	������ B���Q`WE��On�k� ����0��^O�ie��f C��VP��Š6�1��W���!�Ue�ꡚ(?q������c=��x�����|l��jhP��}�y�[��1������;6V*?�#?֮Ү�w	������£ȼ{A]f뺾��򹄽 ��rv������Sm��AL�8�
�+�<\��,� ����*L�7�C�*NS���/<�?��(t�&K��7�ˇF�1�v~=��������r��i�D�٧���4�h5�A���UU�G߳r�a0}���P�%%�>.M�0�
�X$Z���c\�s��~�:��� � ��2�ei��q��B+�L
b��
'B3��y�WhkӦ�� -��w�0��iV3s�ǁ��T�� �kD�����Th���C�6��S�/lw��l��P��~3R�pj���0���J�ϡ����_\{ "������_��ݘ��x�\��6�?�.��
�����Q����>܎��������.��.�.z����*�H��N�y���~���"1�
n��ćT�n��>u�D,�QPf�<�A82%�Gz�a��=�z"�����%5<�ԃ_"=r�N�l4λIj!Ƣ�����u�HH�ьa�q-�%]�Ȓ�K�Q��`��?�Ţ�:�,�Pe�Y���9~�����L�G��̦ۜ�}d��U"�"�Q��\������<"�� ��Dz�����?"@�u�g��e<<o�e��L������P���}�E7�=�yeW �!b�f�N�S�+A�����!��`�'�j��^DC�-�#_9��*D�6({X��F�[�z�B< �쫣�T�{�C�;CN���B?!���SON2��|ܺY����N�_p�3ilg���Y�w��q�V��d�/�Zh0E����c���W6h�,D�#�.=��.�&>BzN;�^���GA҈����엺��e�|{�=0�Ã��7εz|˲vz��7����S���6��䉼䘑zh��%���P��~7v�!�tW�Bf�R�}�����(�<��m���&47n=�׼��,�A:\ݸD�y6����S;Z5i���j9:��M��r7c�����C0���Hg`8!����y���Oߗ�<����U���X�O=U'��Q�y��vR��p�M�U������%J�	���H8�n\B��Vz�~�5��x����Zƣ��k���pDz ���0��`_>�(b�	�c����ֽ��~��� F�QQ��h�R#�^U�g�R�*�bTU�=��M��#i��X��N��j�i_}��>���y������:�q?�B��r��r�F���v�nd�J�~��̳��z=��Au9�aigt8��30�n�P�o���A�|CAr��c������dz,C*�����������k�P�aL��B����9< ��D�G�h�� e,���I��!Y���'��q�5���Y_�m��F�_�hB\�����������܂��Y�R�p����,i
��!����y���Wfﬓ]��((��9P�{�X�8�ш��ۆ��H�J��g��/=�������%	?�s [/���.yC�;�:
��ma���uN ^)q�6_AsU}Z#���B=F�֣�豃M��R=������'z+�|;�0W�=b�N�
������Z���0xͽ�ך`i�P���G�����������1�Wz$R��\����f�ov9��蝂��F.��M���H|�/Zރ%~Ϛ��#=%�"G��+���I���1C�H���)�QL��mW���75��VXA�1�NeO�2��R�j�6��9C���R��1�V���|�m�"��g�=[#�UV���?�;u$�֌��O�1b�)|���S��hsn��N��Q�m?�s����ám�"	�[Hw?���B����%<w�)|�9]�����Y���V^�g���4"�F�qG�e��eɩ:7h��t<#9\7ε5�G�n�a��T�%���j����F��˨���o����1��?6~�����2��k�uV^��
F^˛�@����֗����%Y��Ĕ�A|.U� |5:C���R�O��4�)Ksc]�p�?_�#i�tṝ��Ԭ��1��΅�n�zc��4o�!������T����/(bU[K���3��p��NE܅r
1�|7~�{Md�2=L�\8�=$d(/�(�E��k�)D�R�m~�������uKb2䗥���: m�w�2o����j��q�R3���\��頟�_kq������7�P�d��>7�͝��w��^�ߴ����gpoE�E�/�`B�m����P߃U�E��ᬭHp�{{u���k��:�y����~V��l���
\7</�߶���M��7,*60�m��Y1	��q���[�$�o3�Id]	�h}Lz�����|��-�C���k?�U�M��$f����@�`v��;zw��ho�r��W5�~�5��bx��w�c���)��J}�!��]t��L�)U�nQ-�+=�WNI�w��ۋ+��-־VAӽz�/~7$4�9A��	�ϹC��4c奥wnυf&�˸hڥ��}Stm{[���k��;?���?2�e��%���&�MɪY�_.��+���g�sw��]J$�E� �fX �;��!&��C<��>���'�7[A�W��)+�l��������o��ᩍ3������z�ݵ*P��%�E���%�l�Rl���~v6��߉/ŏ�E��R���Kw�55�5�k���^'� &��"e����# ��i�l2��'1�3�۾�xК�ɲ�+iA��E&Q����� �)�?W����=&�آ����-��Z�C��۴�lG�7)+�b�KF�Y�5�����˙����������7a41^�Fr?����v���_�f�݀�b�Q�D�ԣ�i��*�����^�3�%Y��40I�S���M��W�ag�\`9����~+��U�v��_Z�2?Q�ț�
²�f�)ͨ}�#)�n])�dPCE/������ͯ9F�}s�$Bf#�)͹���q�c4�(<�@{�����xőGGG�V�;ꦮ��Q���C���S�]i嬓���n��爐������>�ɿ��H	��P<�Ż�������4�e�m0M�*�<�ᮐK�Ϊ"�Ō^!=��������s����W7ݘ���I��yêٜW�j��C�i?��/��(py�7��y���	<Y(�x�����I]�n�$n��������L���161r��&6����G�����P{�����V�Έϭ{�x8��?��W��s'G�{J�k�k��0����"��+�|�--��D*���>6CU]z�^M���f\�Nj+�����a�U�x�z�/��_&�(���t|%	���]�5��)�Dњ��SD���J��Τ6y?����讞�]��*Ɖ�c�el6��g4��=�o�C)|�R6���&��+�Ұ)X�������)�v�G&XԹ�&@��y�> ���/��Z��d��g�.����V`�)L�^�)D?��d���Ť����::�%������R�`Uwxh��WP�Du���៲��C��r7�n�zy�Ȏ꡹�ӶNrP�V��j��Z	'�\�`��5��fb\�.]�q(ܕfr2��Ȋ"���xÃ-0�u�����{2Y�p=�P�Ȍ����/K'4��}.��ސY|�I7�`�U����A��{i��bF�[D�3{��F�z�ٜ��V���%��T�+=J�#����^�ŽuX��z��9R�����U���?���31��W�$��������OϷK���	�7X��=�p{����u����5�E$���Zϡ9\b��ڼ�$U��Oȫ!꣍H=N��K�aD�ޖ�l�9�e����:�������K����:�� �U�$T�a�o_��!G%\����mzJ3��X�x�?@RD�
�G#��ɑ�P�A2���}�n�]�+�  ��Z��V�.��uЈ�\�㋈���|��#�]���~<,���������b�J��藋T}�������E{�T]����h�S=+�'���QJ�8$�S����Z����!��1���D��Nj�\�9����$�n�<��z��x�HV����3?%O�{���o�U�21�s�lڱ�*1��Z{=��C]{�3^U�Q��c_�L��B!�Xb��R���w��݉6�T�"Y��Rn�2@����[}�>��E�w+��c�_�HZ$y��`��r�ԥ�'� �M����ذ5���3H��)��ϻ3�I��T&��=���O�ڣ��-�Y!Ds��\��$��T��L�)cb�#{sa.Lj�+Y3���1�74����fo�����Uyc/
�mEr�)ƱiX�ӽ�e��^��<3��O�;���3㶥L
2�պ������D�k�ͺ'~�<"��c�f�N���Y]-"F��(C��4���L��nm� d�='�VޖJ=����]i$����?���D���ڗ��+]-)����r%��՞���,�� q�0�'�c�0�t�j���ș9:I�������rU���^��
�?Z�Dy[5��)T��)7D�v0�n����'k�@.��f���k�M�2���eTs-0��ռyN��C���nm�u1��4D��I
�]�O�m\�"��K��g��e�Ӧ_w����G�SC���^&p�Z���'k�JH7hP��R!�o�3)��K^�8����wtk&�m�7߮W�ti���f��(��or���0��j�����κ��%�O����y6Z���x�5�����`X;�c�l
PYخ�־!�`���%A<�/~Hٵ��r/(@�ƋJ+���-�'�� `�*�Ϊ�*k��7��T�]�_����E�	xB��$"��2��W{*�Ĉ��G�\+0Jx�W���4)<��6w�ٻĽ�,�'.���f]vzz�1����Ķa�[��E�\V�Ȩt��$t��������3���_�0�����.a��qxvV�$7gfӯᮇfs����0�%�P�֑�XJ��H����R����[.�u�0�u#_y� �F7޾�yۃw��z����UV��'|�K�T0P<�Z��e����&fT7-�^�}O�U�$�0E&�gK�1m�����ʨ'c)��:oMPt)Ƀ�Ȟ\G��Y���sL�̄��r�z�t��=�2;�������3�`�sp��s�y�h�b�:� �85`ְ�� �6��[���W)�'�k؄)n�m��"�y?��w���	�<)Md�ĔgH�N�
s"g�L�����K��F���,���Ml̵�ԵF���� �U��H���`ֻ\�`�Z���]o,�g�;�H�p��\�`Ɵ��GM�T�҅:�2��d�n�D��5޴W/\�P��]U[�]= ��&-�-���S`��^t�"���Qr�r���ֲh*��w�Z�>�����py�\����'(��{i��KӒ,�-)ʉ.�(�"��e�T������]���\�;�ަ��:���n��'&�e��)�#�;���{Y'�@��QY��K�ڠ�}+��!NW#��r�ۑO�q�%�]Z�!G�t_���u'��B�� ���}L�??i���i�����;��/U���������=�ݧZcnڈ><s�<�P	Cw�#/��K��qO�\����Z�_\nY�	�P�!q�Ф�,���囑$�v눁����A繘JD��=j1�sX��}9]���'M��u��^�A����Yp�D��������O�ԯq����̚^�z��`u ����il3J��[Q�D��^}��s���ղ�A[^���6��yd�KFv��~v���i�-�@��r>:�:cܠJg���&o&
d��ȌU�L�z�|?U���u������e�?��t�n�r+hu����6{ZZY���0D�A4�+6�2�"�����W��j�7����q�#��Y�m܉.k&YЙ�2�I��A� ~�ҡ�v�9z9]^#�v�ݒ5/��[ ��z�b�ǀ���7ʯ��ak�-a]z2��_�/\����Y1�t���U�F�{ǆ���x!�尨w&�k� ��NL�іш�Z�7URZ���I�Ѝ����8��X);��@nNJ���Fd7�
g�6���Tb������3Q�7��)�������FG�s4FՎ����*#C��סZ�0�u��3h���ȥ$��70j����gc��W�CVn)�(��]�����0Ʒ w=?�ݟH�h�5����RuTJ��}?
�:�e�*�4t@���J�7�U��b�q>���i
[a�G��~������B�J+N�5��,<~zn|�J�X�(6ps����W ��\򪵘�Q\.#n��1��|2�X0���뜪�IHa)�I�H�U�i��}�kn6J������LFk�3�GLc�����J�����X�~ڇ�Ç{3�\��m��Uq��>N>�T���ż��NN��C{��u��9�̝G�v32����,6�\m"U�O�:�{7u���*��%�;���d��Z�o�K�c�fo������ >,����e���)����t��� ��RK5�=b��"�
Z|/�6�~ �gx��]�%�����)�$ݻ���_�.N���ƿ~����٫ix�&�#J�T���p������2|A4�T�����-�cf�����1�s�g1��l2����_�����ڠ���1�1Ħc�r����̜`1�0P�EJ�j�x}�?e�F���k)��4��x��5�����*�Z���ܦ�v,�&K���ϩ��Z�h*���'6�[2�2x�QA�h��u̻����Bx'���o�6��a�0�.y�zrkb�ˮ�]s��OvΙK	N1c��)�����4]+��Ģ�71��~����E=���E}�57<_�6[�F����u'���w�����
2�'��K�񮄁���r�gs!aLJ{;v�S.j� UaR:�"�W&bl�qy�i��<� ��WL��ظ�G�>�+�qn9 �Ƣ��M4�{�{=z�}��c1K��|���ȃMy۵e2:�d�B�����O��s�1}�w��Iye.��g�ig�Y����R]�- �K��=����krb�I������a��ɛ�����|� ;=��%	��&�L��}�'n�,���wV�>>�$�}gώ/���z0��bR,!�g#�̯�Y�p��Ϋo"`�s�G%<."=~Ա���k0�/#&�dk�DP��ES�R��!��ӗ���p�\�C�E�s���̲S��~����ni^�N:��!��Ù'�<�ԝd���9N+�!i�Trç>�<�� z���}�B�{��E ��pn��H�2��K�op]���`���K�d��෹@ʂ�\��n�|�g���
�nK�������L)(\&������I7G��	��1`��)�X	�d�(Ο-CE@{!�-����_[�kޏ��9YQ���X��x[�$�R�XΥ��I����R�������!��1a#��O�u���q���ℎ���T�U٧��s��#�'�'�����T���?�dj��L���卲��ڀ���9�U�CK˭�λvైr�|k7��[j���P)�;��ocf�,ǯ�P��WYr�G&aXE%�{�Ѡ9�QL�|g�F�#��#��"�����/��X��"4T�7k2�$�i����Ny$�����Y�G4�}g:�Ͽ{�<2���ϳU�sRa6O��[n"ަ�;�{� ��~r�]'6�c�����4�N����*^A97��M�C���M�suf�����;R1���N�w�F�3����v����'�.q&@L����^ӝ�(/��[o4Y�:�YKm�<����:��#�Wu푻	U��b�$��_/�	���ͻ��g�|�M�������DI�:�/�f�)i+9��iLxF-J'� ���b�CO��K?���5�:<spx1����ȫu$����F6�!�0���B|a��K�J�nsy>Y浾g@�(����UU��)h2  *���F�?Z�K,0�H�7� ��C>�4b<�f����!��׬@M���gD�|N'*�Ҡ���#[��������t��$���F� �"�~NQ���X���OD',,(J�����2�����UN��#^�/I�o���0���!،��˹���tz=�U����޷��M%�_:�N]��T-[���j�usH���߬������Wp�0��V��l�/�t�ĺ�ˋC��|�jz+�B�PK   �cW�����8 �I /   images/31d687a0-e383-4fc9-9100-a6b790c355a8.png���7����D�D��D��	�k�{�u�!D�-z�h���3��� �`�2�6��w���'\�~�΃s�s�{���k�=U�GL����(�Ք������H����/���!qQR�SWR����rtqw��*������#|MDN���N�X�M���#*�(j���d��z-r�
�Տ#�,��!@P)�zO���\N������-rI���"����{�ȥw���
���j�St����?����-��KV�� �O�w?�Prd��:��z;y?�f/}�!�4&"�%%i,�%'_5cdx��9`H'(x�&(�.�J���h���c�����Y9>'�d{kꮞ���d$,�x H!';	�ї�}Գ"�`�Q��l�h�h�hF��yyU�=<|<<ueE� �#�S��I�z���uut����C��<����ԋ'�{�@#b��Z�p��Qq����B�s���\�UhW����+1���s�����G\�DE`/k''sB'�Bέp-F;���������?������?�?�DW�{�H����?q�Q���E�������@z�"��iuu~�Ԕqf��!�G�C�f�¨��"G�*ٍ�@  d&
��� ��:V^^���5�c���$d)��4���Ǯ���(�Kuh�ּ��s�1�l����}���l�^GM��X�媄v��� w�u����A��c�W6IB�`l�
����됭����@��!D���C��_�� ʹ w����heeX�16.Kd�`���ް���p�����Y����/\�l���D���oR-�v�����n�UO���*��X�#vܭ�(� \ɥ�b��X_�/�ǃ��ސ����wm�'��
%�� Pc�kD��K�Z8�L�{�xK���TA�Yhy8Eq}qSr�vX�Ⱥ&}y���M<���o�����=����$�V����@08���Jw�a�-g)D�Ep� �J$e{|������к�yբ� /;�M'�@�ATx�$��J�Ww�(���:X��T����+ޑr��xa-R��4t^#s������F�ӆ���>%}�mMkP�p�|w}�ݟ�ӯ�|H���U"�
��iQPa(����sQlvaW�u�� #���U��11�iDêۊy����L�]����ς�w�j���U;���:{�U�nA. ED�@7�쓌���?�NR#]�=�_����-bKB��WD�2���2�-�Sx��ۻ�*Ȯ {�1�k�nHׇ��W�v9
o�f61�聙K��e �bn�nvxX=�æ|Uy\���_�MҭH@ DD�3byx�O�hBT���C#{U�S|����̋����f��ZL������{ҋ�s�DE���������:U�"X����04��M`.i�Z��|�_Sb{A/��i\{8s��QM��:åCJ��T��I���x~�2(��l�E��'E��������ದ:�4U�y���ޱ#����BK���1��1�,{%�?H�k�#;�b���p�	g��x~A�T񢡓Z����ݹȻI� m^�lsa\[�-ιN@ԩx�{Qƀ.>X5��_2sⓟ���MU�6޼���c ���e?�	��z��O�g$����f^�s�C��R~��28E����B�����=��;Lt�G�>��M�l��;�uI`0B�����/�W�~S���$�)���5X>�����!J�%d��]��K��!��ՈV82=`�ז� �\�^UѪl���ۻfw��wtd'�2&�R㐽�1Z��3v��U���
@�n���]p���>�������j�&���F����Ǧ���O�>�������TJD˯�[�6*)�O���'QV֍�27�д�)QR(������݀-��8�s�1s؉Xq�9	�j9 ���#�ww�b�8�	�_l"؞�4.�~��d���Zt�X�����:�&�����Q?�>b�u�bV#`8kl��KR�q���Z|�֒~���f��=������!�3�'-�ӡC)��D<jo�����ǵ�0�������[Ug��7�;|��w��L����c�a�dd�܏E܇{9�9�Y��}B��7fF�z�YY�O�y��Ԟл���U)d`��O=L�:��Y��b���G�L��xN�K�������)������ӹ5�n��V����30�i�����2����J�%�J�Y$�rjq����z����ɳm����9ttt�}��x�i/x��KE֣{aR����3���r���h�*Xު�M��&uE@�V�iD\�HѾ.�܁Qfc}��.��O`)k����n�I-t��p@�pE�xW��)�Y|[X����ѭ,�ꔨk0߷�>$$t8���	�����m:����Ί��IA��?�"��3��h��ٶ�&�^-��k�����AS^�s{�������]�9H{����s��gӅ~�����W��[
�[Z��[I��;�h����#�]�m�Ϗ�Ԙ$v���Cs�T�^��gh��-��͟�R%�$��&	���i3�9�d��_l�:GH��6���Ȁw7���ݯ3���˷ĝ�����+p³�⫿&���S@Ѝ�H����M��$yЏ���v�1�����wM 0X��j��ʁk2�y�t�����D���	����h[�b?W�n�QNPZ�2�c���L�L]�R[8ͦW��Fd�4���6��^t"�xt��[ݘ���~��1�*���7C4�N�e����Vx�n��4{�ܩ���*�Q�(#�Θ� �t�߯k�z7��c:p�v|���u�e�ӛ3����˲^���
Q��AW�e�@~
"��	��Q�Y^����m�ER�Q�S�(������.������[�ыO=���7]H��吊�I�n��y��a6+��J�lٺ;�eZpCfS���X\NR2dg������P�B�Lh��㪫֚���R>}68�����#��~�t�U飘���.��0,VV�%�o��5�X��6ʂ�t���yd:w��s`����v�^r\�`��VQ�ƴJP��;�_`s�X���fyF����ׂ��6���C�Km��:�����۷���}�#����ǒ��G�YM����r^�<�I<&�oþn���4Y▏��r�|�����l~�\��"[Ĥ���.>0F��I�έ��p[�j=|Jl�l���g^��j�"�-+�Tm�Ŷ
�� ������TQr�e�����kH�+�-�[�����=A������H���g%s\q����8���[����\�v����Wx_��C0F���(���_U~QKQz�|S$&f���N����ܥY�5�ǻ����Ԍm���f#7���t�����K�����~�&�
^�]���ZY� /ɀ����
V�h��B:bguj��L�A�>���Ƀ&���_�ߍ�)U=�11���Z��%���)K`����I'g۹�w�]/���V2� ��
,�v3L|�d�G{U�S�p��8�����U9ܹ�9�Q)㌪��D�R�L��@b90�"ڹ�(�GV�y�_x�l�۹k�#(���8�㵃3��W�l�P���MS�^��7�<D����ijsz^o�L,��!����>�L�kh��S�x�0�2ROE���V��l���@�%�%��G~s%q�D����p���1�قD�t�V��(3�ɛ��_�<e����!7e�I�Sq�=�c��K����`)����d�g����҉��g8f+��Y�LqLK��%�))���U��� �"���[=?m���q������e��a씏ceמ��8V���T7�Y����#��?�3>NX�>��l���D�$qg�S���Ͱ�R`xܣ	�Ds����A���-�E�7j=�h,�����U׉*ї�C�]k�	���U88�gtz%ojZ��GY�U>\:2H,2�0�y:�+���H�`�������)Y����Ta��3af��	��%��������kau�<u7��K��R�`�,��94�8��xD�p�\6�-�۠��2�l����f��p���n�B��šE����e��Ĳ���&D�p��w�Ȫ&#A���t�p���p( :t�x�M���������¨�t�g1!H��f ��v4&�0��:pE����:Gi��[i��2��Kխ+T%o�6��ʒwm��t�~m~;*�ټy3�QY;���O��Ή%ڤDl-S�|BT#��c�SV=�&Ͻ��H D��������Q	�B{�+k�Kă����M�G��SP4�Y��+�U���Y�dj���hRR��� ����՝0}�����P�
m�����eP���DC~k�WPv�|��Hϓ��]G�/�@�%�ȯj��q��?�EO�,nv�j��K���㮈��#w-r�o����q=,�P����������Tf��eI�-
����;R��6�F�ƙ�޶�,�����\`�����	�s#��%F>��j���
�ඞdٻ�e�w�m������5q�{T!�" �X�����s�v�*tc��6b�m<{0���/����1X�y�_f|�7�Z���:�&S���*g$���_<rCe���n]PQV���VfT����'7ݫO�{mݭ^�g˪�y� CEіӣ�-�J�WU�)��� �ŎQ�Vw���c�q��c��F���#,̝Gs���F��#���tQ�P��GW1��"�`��9(�3Yq���2n���u	���]�� .zto8JΝ������O������=J������^ƒ�ÏW�7l�F�٫jT�H1U�[������Zu建��~T���V �݋H	�WbX�B�شa=^R�˙{βj�y�KE�]�pi�����{XC�S�V_T1n.���#~o�$հ؅D"��q��u�$)I�).NVM��fV�Ds���r%6��q�✧i|��Dkgn�Ov�%�r����zx������$�O�<<2��q7��`1������:剹C��J�LC�b�b2��]���:�1	��"���7���u����ɐ��Z�9���
=W➖dvK����0��x�Xrr�p�c����Sǲ�qYYH�7��p�
����5�n��3:m�Uh"�S�T��h��C�M3I7�9r��,�`�Z�UNEҹH�1�]��������K�_UPB5՚w��n||�Vڷ���e�?u�hXᆮE������P:�Ϗ�%���d۾%��
��,u4��$_W)0�O`�u}�G��p}��$��s��Q��T���x�X8�/Ç囖&��?�����׭�N�4Yb4�K�q	�N�"M(=&�����E���ݶ������WT�����E���؊��A�I����L	nB-�)�~����Fx���Z)0m���R�؊i��K�zc-�6�>�~f@�5zHՅ���Te��0�ٸr<���^��^Qq>
�N=��h�զ�ǉ�p)!��z�(@NI~��Q���Ru��t�Z۬l��}&:�P�a�7<d+�t� �Q�E��Z�A��SX�un[j��6B?�"�'"��s��:sw�������0�w��I)����������,�	�wD7U�||!\��I�'}%���g{0���}-(��MDH������������t��I�$�e�á A `_׭�,��=������UT䠑��͙m��+6r� #��*�0�t(�=|�.`���$�:< �>n�3*r]�.�?
˓���u=�@<�1�bd�ʿ���D�L:��6�́�*��d;�<h{�=��]~w?���]��l�w��34���X2���(���f��W{�@&CY-p���b�`A���*��_񚬟�_�>��g�VG�	ӓk-�i��c���eG�ꠙ�9�!��2���N�
yR�z����?'��>�̹_��po���נ��]]�㼭Ǎ��8�
�H�9��� �8 ?�uL��`�>�,��,VQyMt�a�����kx�i��ql������*����@��̄���a�x����݈����C �M����.$4��K#[,���|������U�(���2�}��r`�F��(Μ�n�3��y�\7Wo��5��mv-w�)!�Qk�R�5�G�ݚ�����@59�+�r�������=��C�LN߇C%xjʅ�8�)�?�M�Gǲ�G$���Q���:��,�*+�q�I��iC��[;?�z.�K�?\"������d��n{�o���m��q��8ŠW�0$��P�����Z�*|M-SW�����9�?D�/$��V>g�G��9���J��0/}���,�9��ϠS����b��Z�mH��}2��Cz�Y��?�G��U^p���e��3�[���=36<7��?���K���c0/�F�5-�V�$��ԙ�r�(7��;"��;�G��N�s�`�2<v�A�o�޶fWm����Ѿ>�#��qsj]�������ě��׏��[SL͹2)~�nEGg�7��s��
\��0)z�S�R;j!��A<Y��!��4�X���B";�n���](x�m<9�/<J�>J]�����.,"���&�Zm��/�%2���EG�K�W�$���9!�"4ز��
vѷ�Ȥ��|%$�����n��)藧�vM��<�#t�Q[.��V�]M��˳J��>5��O[0�~_�*��o���M�=�m���/��n���h���\�J:��~P��PԟtS��B=](�$.��+<~.�>>0��Ì���r
ڃg[�L��34�:��У��e����4|�]�!���~��Nxd�%���L�G-O�O
x�=Wgɥ�M��s���a?+ʈ���ĺv�&�!{A�=�,-�+煮B���	���Ŷݯ�_wc'+�o��R�~�fݒA�$���� �����/z���d�[ЃXh��0BL	m��H�hk��|��w�];23Cn�@�P��o"�:)�:!��,��`���V8<��P�'?;�y��<88�d_
�%��W�o��[M!.�qS�Ǣ0J�����to��4�	�2I8��<)kY���+B
�%6�3fk�w�WO.�_��p��߯�;c�_Xל�r����ʪ3������Z�çw�`超>";��6j�ʵ34�F�si"0��nAA�+���v���ʜh���\��>����Ϥ4����^�\�~K��y��``��p�������PƋ���btt����l�E��r�,嗝 ��i{/���R�ԃ��O
Mp�I��5�y޳'�#T)�"g�n�uv�5�)��a��C�?7�Ƌm�y̄�'�T`E ��H���w GlX��슩f[}�桦�4�dڷ"����&ߙ�E�C���DB�ښ�+A�_��V��AD�VR�� x���Q�Fs?����$��*:�
��z��s�Z{�E��Xu4���� <u�&W5�!�g�GӴdd~�nۇTlK����}ź�,�.gҙloyV�lr:��Y�Q�h�ά�ö�x�G7x{ ^V���9�����#'(�ތ����J*a��\��C�>)"����X}��h�b~:��������*�Ֆ�	pfh}�`��Ώ�ˠ�1X��v�A�n��*���N�a����>����[%睽��4�*Q�;��y����=�1��yDس
�$0񩛠��VEIzI$,���$���C�MIVv���G��Sw����&/���Fܕ��/��'��3�͗$k�Qȱ7���aO����s´��P��t_��K��fu���E5k��-�sKu��dX��t���)���f|_��V��$��ۣ˱�og�uՊÌ��V�{�k7G�va��E�w����篘!ѐo%�)��0�8������x���m\�%�)�b2]�{�%t���������{�������l��ߍ��6N������Ko���������\����v0���K�;��2�<���ߜf@-�2����u)�XT��{�*�}��k1���b���#��73<l��i�t�{B�Ɗ��B_�HJɀ����NE:vs�Cr>S��bYS�_1��2����Rƛ$w�2VL�2��G����>�к��.:�s1�����x9k���%�#�S�Y�� ���GG�s�dQ��ȣPT�:%�LYL{oɎI��U��1�yTZ�@�Atc3�G�-��9E�Zw����Kd�wkJ���UY��4F�O]sK�ר�ef���ο�-���-�%p�RY�얮��Mu��\�\lJ��p����P�bhFh����cK-d׌�6������+=�e*ߑ꿣��֚_�����v 4&�����|�5�{��'P�7���E�@@k��d����߳F�	/aӋ�Z�%�a�,�<��_rF���;��������
v:��.��f<l!#T�N�(�M�T�Z��f�q 
���e쳠�c��h8q��p;����"�����s��`�*R�'_�s���?JP�x���d������[\
@�$�����4E=�M- ��9������kU�]�M�V��
��v�@��Gu#^�b����]���|
��>}��af?���
��g��"^=֨:|4�kY[@]@ǭ����<ld��HPz�ό��zh�b����+�[;�?� M��gm�`񇸸)�S���DL]z��f�����x��x��U#��R����R�j?�2�3�8����h��4��Hn���<����^��Ͳ�P�p3�.�޴�X���3kA&��FdD����2�P3_T���R�E�<����/q��<��O�n|�%cwc�DQ)4�`�O��i'Q�ҦTX6���^\�3�;
&�B��47Gy�n��^3A�	��*��)��ݦ�o�x���&g���.��3���y��}^��R�33�0���aŔ��7�ݶ������r8�R5�jױD�6��X���je�W�y+�2��b(+l,��~/�!��!�&�)����oB`��[�g��Ȁv�M"U |�%����șX�$���~�}������6��lB�b{��Ŗ��Z~�0���}��ު��U��	Ct�w�z$ c��e'���*��B�n{R�z�R�]���I]-�"�j�7�S�#�BNt��H_`>�A6�8yR���8���t��;9X9h��+�|�q�/�4u�M��~��mf�ȣtF���k>�>�,�LeM���_���灶%/�� �����(O�
�tqS��5�R��$�>��n�c4<��N�����O���G�Ց��e�-�Ԣ7���E��������F��7hvu�o*L���(9ϖ�\F����{�e[Ϝ
�N�C�{{j�T���-)1_)�ٲ�j���n�߽[��G�@h���(���,�t�Z��������������ce��q��8�	�S�z�**k� @��Eg�"��-��/澝nRw:�-$zr$s3��ӓ���ύ�.Pz��Z��爫�R��o��l;�R@ݿ��:[
�d=�z *��`Rm02m��	Z%w�����T�paw��m�h}Gر>7����ۋ8�h�/N���J��"�g?ُW�x�_oQ�ݨ���@�o=����~V��l���6��QB�nZZ�ku���ab Z�^{�t_@�*��Cy�>ޏ�k��Y:�+g����M��f��,ox�h��c�?��	�O�����|B����II��q������OH�ꑲ�_����ǹY)�F��CD����aGt闅� ��*3c�������o�-�DA�>���.c-�$VD��Ry���
��[ټY.��Z�^�Ye������{�b��B*V6�*K-?:���C�먟sq�>���̺v�l�ev5��M��g��裃wT;�GH�(�5/���TV߀2~�A��J%/��Um�(!h����XY^
�n'ܦ8V�D�t�N��4V���e����O���_RF���G�_aj%g�	#�fs�V�pψ���_MV}�F�3��?Z.��g�4�?|5j�,Ș�Q���'�;*Ry�[1v������v;�}L�f�[3�B�K%�GSt�~X�K+1��6N��:#J�KT�������(sUF�3���F��� ��y�qO<}D#-bF�Υg$/�³K��9�v�#;Y�����?èF3�u�~'�r;ו;}N9��� P ����T9��{�*�yF�[�2�9��+Hw��k�V8�p��QXd�m�^sIv
�4�����_�|f橅!W�-�;1�@�X4����Ʒ�"���"��<�]"T��/�ßM�T�}�"*���:Tώ���.S#m� �zt��e,S���*��vX>wL��{�iכ�f"Gh��V�PCEGl����3#�Q��[��^��~T��c�6�x��i�֩z����PYy��D��3���A%�(J���?�V�˖% �a�}S롁;jX�M��;e0N#�L��`gKQ�@�����!#�W�:�і�Nl�[~�8�M��x���ϝ4	8�{�:]��rsڿW�v�R�.�,s- ��5�%�&
�ssZW�u�
w�_-f�� _J����'-̠��T���A�o@��'O���kS6E�%�ȗ�2�=6Ui�kW$:��% ����L�o
,A|^]��,������C2-�<�T�k��dV{Yd��Ɣ��u�go�&Ӓׇ�_���4��`��.�LJ���i~�*n�[�����t� @�Re���?��wݸ*��i�T-��ws"9�9]h?Y�L��-��C7�	/:��[�����sw:WO��u�vt����p��T�ѻ`��g0y�����b�Ƚ���ȩ�dU(�{vX��h�#���(z$��0ןe�9�Ӵ^�t�D�����}}�<�֚=(��/���I�����Ȇ*��	�&ٻ�F�:O�o��\��Yq��Mܨ��>0-��:�N�a�9t���%{9�U�0�W��O�bsV?YU��Y�j��HA�"��}檂�^��4�
q��QBF�m��&	�͕,�Q�.�#`�����J���2�O�̧~�-��ȁ��T=��5���W$�D�ب��A�`~7�8���5�\gd�X��%�����<(��=*a��y�P�
+�)c19�c��J�WN'	1	A�fj��[E���u�Qn�>w�;fS��n�$��Q�坧�'=��z��ք/`������%[~��}�:q)�r�D��Z��6�N�XR��tPw�G���3:�m��d.h.��g��
���2��!OR(cf�uw�*��\���c��1��d:)�Z�a� ���W<1_��9f�*(��q�J�<���/�/�W��$�$��yZ���ο1e'���Z��6;%�2#q:���:�n�ɂ\�`p	Cn7������,����ãl�JO�2��=���łF�m�{D�T?^Q=�*�Z���!Y����rD�w;0J�<��<G��pYaR#�{qq7�G�7��~�o�w6p��5mËb�q�1�0��a+�zI�Yv������LGE���P�{ySԳ~����j��Y���j�K�f���-��=��U�(Dt(�^ߞb������i0���uk���ڴƩC�v���H�Mᅗ'4}?�x�u9V�;W.ʟ���`��Ӈ����"�a���K���8��X��v!���Z�eۿ]b��^?�"�	 ��B�^�̅�Ҧ�ž뚈3uq�}Yj ��J �!�Ȏ�Eg f�.�w���<H߰2��	���P�h����YJ=qx]ӂ��m�ڂv�4��+ڪTIU	6`����&[�T���u�ؕt1n�ě{f����5�No����Fc������A�i�ݧ �'��j��^�9���9I�+ƝR}v�4Bb/%@�^�!���f�KK� ����Ft�c��"y������D�>}���Z"�����Fv�V���JO��F��������44����W�F=���	��-�X g�e�<�$E�o�7��y�m�<Ga5��!�vz���wL C1XM����n�Fc�o�KZxѣ[�y6k�-P31g��r�}d�ek��r�#�5X�i$)���EuTW��nMZ���$�}�L�{��W��DD~�PP���r�!7���/*����L���0�!���M7�%ѥ���O�.콢��a,��ѬǛ���b��%����N�kx�5y����1n2��Z�w�>��İ?�b�C�8���i��,Xٖ�=������O	�H�*q5U�z�萌�-!��\��or2d���t+5��s��\H�.&R���ӆ����,&���M����l���NK������t;G�w���V�C������Wv�"#{_C��ֆ�f�G��n��X�陔�l8�����]��8�0�axE�,/ǁ�V��X��n�6�Zʨ��8F��\ �nW��������Wę�Bn�2$�r^$�e����j,ؒP\q%u[�#�q���*<&-������W��VVf�Ul�#.�m���"k���yR�Ѓ�݁@P��Z����#�}J7%�a"'�O-���[�X�a"5����}�F֑��c����1g�o� Β���N�Kըl�]]%�'�"���A�H��sr\!�f4Q�u �	���;�K�18�ݖs�����V7qΧ>�K#�r� � ���0���ag��y�cʖ��[��Ul��\Q�iP{��L�#x�xMv�= �e�F̘�R���O������ve#��mJ�.p3GMR�q�<4d�(��C�͂�<�Z������ t��<z�����������~��O�r����?����i�C�m'���j0}��A0��d�Ǚ8>��A$�Zͱ�@屰��4��n-F>�ޖ��%�(��2K �O����8�w\�MZ{��T�8��D�(�1�������6}$ ���=S�������Ji�+���8Լ)"LWv��U��l�"%��Sf,e�{me>�3�h�����M9Q�X�ȭ4�G�?�5l{���������S��_c��ԇ��H��|
zBl�Rc�x�q�Y���P��mE���1՜��*�4>;���4���iM|�MCIlz��D!Rz4��Fh/�/�����f�mʭ�/x�!�ȏ�w��zCt������E��]�̫��˞7��n?�A������V`Q����9Y���0�T���6H�}��K�=��8�6�����J��L�m��|z9�9Cj���{V�͓W��������\�z�X�tt�.�z_����
�R���k^̰�X��3$K^6�X�C���*ο�t��ʿ�*�:3��35_=p�Q�L H�ŗ�X�ҷE�ח����7&g�A"��A�-IΪ3�eB(��'�-����+�\0����� s��"���Z�ͣ�N7���s�Ǌ5]��(<�{��_���{欁��P0�O������J��^G6Ǚ?�ƥ��T���K����o�������I���W.�"!��P	b�2��zr�-I�f���8_�s�d��K���a�"�`�G�vM��͔�J� ��r:6M��*����̪�S9zuf�7;0�W�B�񹏭�žvD�ؒԄ�%ߛh��A(�R��=�-t�3[¥[1ڸ�����vb;ʌ|]:9-��K�n���"�1��[��� ?ѺDQ��h���\7%�����DČ*{��>�x6�3;��*�!6Bu�[ufZ�d�w��߮��7�m5��T��m����T������pܨ�5O��?K!�B�y�b 葽����x���4��@�V(����.LoK8Yl�p�Ö>	ƿ^/d�n�e�z�lD��b��=9��"���u ��74�Oa(F~}�66����nL��9D�� Y�4��g�}h$�����@��-+�e�x�P.���!��^��^�x��������=�A�U��{yX��ja5Y�w"�f+[�E�bu�}:�b��V��/%VY��\����^΂�;giq���ҕ\hΑͦPv����g������GG��?3čH��r�*��MS�٫����@�5��_n)RF?5H�t���t@$��5l��v���o�`'���]�yJ�C�19[�/-�;^�M�x`�C�l2Lwf�R+��eA$�͛�`Z�g��/|@}�����C���a���f�"�y3
�Tna�g�y�����؊���'��:6vվth�y����wH��ۗp�����dj^�m�XJ��BB�rF�:m�S���#�F{0}���q���<�a �/Gϐ�&��dA<�xA�����&�8�D�t�+���5�����ՙ�B�ON��'@s���v�O~��g�xEx�����]��w_�P{Gϑ9#W�i��w��؏�I}ø�I�%q&9��FL��𰝲��E�n�/�g�аPU\>n���6����[���W9��&��#6�����7����r�;�����e۬�}�@���\H��+�k�puW��4�!����i��ߗ���R+)Qf\<����,��Pa|�����@{՟c��k�t�oۈ��v���4b���G�ɣ�:S�L����V�����
���+���r^m*��&7r�zCc�	s?C[[0�a9��$��P��vE�l�6��]���k܄M�j7Ý���e��iKͺ�?R�B��̒�����j^�`�a�Q!���t`�����e��[����l�9�|�����KO����D|�r�><Oe*�j�4ry��B�h���������wm������m�Gͼ1a-���E-ñ0�������]ˎȴ�(�>Z��Z�5��]m�u���}��]��qh��|�k�?&]��g����(��孓��p�C�Mn�.�?���TYWq��&�r��g�
I[�r]~�G���ɽǷ��=u
�!F�0k5äL��#��<��*.Gq�"�2�1l��V�O �<sZs�*a��0����'�(+��Z��/�#6����7~Te��Y�#�N��S%�^ra���Q�N�i�nBL; �j��U~�)��ث�n2Ҵ�e�]����I�=��$2�|M�W�90n��xD�p�C�J4�L����"%h/���"�?p�u1�{����J�;��(���<e��ϒ�b�m(���S�7�XЪm�^��ur`<(���(T~T�֘vDp�I7��.A�hx�˖�p��X��ۢ�,�T3�Կ�������3����v�9��8��^�y��t��%r��/!���t�{]<;h�]j�Q�jo ��t�R�z�4��xlh�1_��36����ԗ�>���8��ATv=c�
呿P?ۊ�&���Z|M�S�9:KcY�o��|�!�ĿRņz��+s���d����Z���g�?M��7�@���b9���]��$�䑌�)���x�{��%>�$j[�f�Ϝt�7���X+W�O�m3�x"Q���9u�p�|�$<�������-a�'���D��~r��on�4.tʫi���JOBZ����-]�N�� �&D��^�9`)[�� HB�~����%7��n��V!*U@�������l�"yz�~?��*���}mE�
�̺a��8��f[ha�q�6�$Oi�d��A&��`�w,�v����.^�d���w�Л�o��"�n�dҼ�nf6�K�#R�pS�����r����S*�"�@�Հ�4�3���� `�7��$$���)@�|hl��J�:��uGa;����-���z6�n���{���;��	�g�*�'�c�b���	T��Z�S&�:�?d%Tlj�'�'�?�	���.n?��e7��H��HWLĳ%��6#��#�-i��#dʆ��|����Ky3���q�(!�,wb���["ۋn��ٗN=f8A�G��Ǉ����<��յ��?��;mf/�,ī��f�yD;J.NV�3P�Up���)�Z+	h��kE�x�K%-DЗ��.��ڥ|b�����Bc�4�Ҏ��:uiY=����n�\��tZ$�ʽ�4s<��k"8;r�&ة�k1��gX�KD�{�d�#�@b�hG싴�GiE3�C��b<�e��{��vbŃ3 ����6v�eU!�w��T��,�Q�J��_Dɋg�QJ�A�i%��n��Y����C�G�Ԏ 'Zb�7��_���Zl׍
�Gɦ`��oa("������v9�6?˔!���é�$#w�39!�#kǾݪ:a�)�B���{����(,�u�L�[aQ2�����+�҉=��|,�K�-r��@�򡼢�T�J��Ik��z�����խ�O�K���L���	��#F[J�yP!_u)�s���t��d북X����B�n_��%�����QG_㾺s�d�����x��^46�k�+o=��N������>^�,�5��.�s�wk�>��;Ъm����ܮo�w����a�m���܆���t��S�Կ�l4j��D�� �3��Z\Bw�q/� �q�j|
�J"KV��_�$��H)ND�sXkrc�r},��e$#�I���d�|����t��_�H���6F�~�ʆG���:��Ag̯J4��w{�갂R@X;��x�3k��Do�0�a�$rrwf���TG�$���pU�F:H�#.9�P�!c�o��C55�ź�A�=
yj�2R���	�á�lȒ�,
	��
���.�=N��&�a<r8�ƾ�-�D.E{�S��#���"gL����3{%���7���sYY~���U�ׁ�1q�!����־�H� �*�8��׼�3�@��f������1��N�Ző��a�J�s&����Aj?��nr��v;���dpV�������������?�2�i=d�/W�M��H����04ѓu�B։#_��9m��;Hl�6��=��;WΥ�6����CQ��Ork��ŵ�8>hk]\��t�� �"|�3������k��HL=��`,߫����@�=�&�!�*�������ԤA:s��@?<p�ZZ��b���V�Ps���8��k0�WY4���DqXca�Z)#�8e/}��~X�P,.�%ޤ5�:�Zdy?���iY Q<�#i��� �Hb��5_(�F.��Y��pJL�Q蕴�F%׋��۝��r){�NK[Y]B�g>���n[�:#���#���i��U�bOP?����6�0�ylQ:'��_���u��<�پ�IP������D� j��y#����A2#�!/+k+���v�}�^������F�H�ݥ���Y�Y����`q� ��h�a�R�G��ym��m�F;����ae����׬5Z��4֘Av=�i��j`p�ϰ�v�������>����r�¿�h��b���'e0�F��Ӟ�	�F{����![KD^���&��"T�)FD#8{�� ��]�Z΅���A1RU(�l+*�"O��/��C�p�-���I;���y�bwm��<!!���P�qX3�;�Z�+rOP�Fk�M��R$51�4��KSB;(k!���u���jzȲ#�hS�'�/�Lr�m����o��D���m:�PT�~� �{��d���'�*��b,�-��X׀d7������FMׁ�5��Q��:��IY��ނ�5	���} �LK�{���;�%�U3��RWd�}׿���{spO�K�����;�	�o�]��q�7{1���1��w�fSvI�^Ľw��Sn�_���i��3d��5e���âs�i��Ak�|�{H��'�p]3>�����B�6��p�zz��L��+d�S��V���`@�[�v�8��0��3�5�h�t#ǏN���0�c#=��#�*>׈�C`}�ѓ�2a��A��j���2{me1�ߺ��o�F�!�i�=<���D�:�q�bh�t|,���2-u�Ř�1����DH�k��"���<�G���*�H	�T.� �9�ٍC��A��{������Y���=(�Z�d:���>^gz�s��[i�܎����i(PD}l�:}�wX�d��DcoXsچ٤=��`�L���JD�A+��w"�gA��wR��l���V*�X�y�h�D;�L�*�0��)L�P�� ����������j��7��/��/�g�y&F;6�ܮt���P&�]~���|��X𖦙7�m�����|x�: ~��>�����U
����a��=�U�e��@2�|�
{������������޷�n�{a�Clo����l؇�ch�u�d�4�F�UcP1�\|� o������eh�!&���q�����B��en�`XC�m�uy�{�+�n��FT�Β�����q�S���8!@�v�2*�;�*X�$6F�zlL��(�u����*��樓#�b*�1JoB���V��1���3�Y�o#'1���Z,l���y��-r�U���:YÙsj�0U"�0k��;�ZD�*p�F��	�>J�UƯ��.eX�#�7��� 4�?�4O:rd:�H�7/P�9�F�)9���L�z���p�HW:}����E�Xt��N�9��kF�B��`�?V9��Q�,��&N�'��4����^�LC�v�*Ñ��_��/�O�3�O���q�Ȳ"@U	�tr�`�^�C����V��_1�U5GԩۗF�k��KvԽ��+U��s
-��v'@ bv�zM�GK@#�g�ڿ}�n��m]����7�Ҿ��,��}��5����6���Y22�
�[x�.�rU��L��}�H���?��_x?����dz���r�Y�=88N����u�������8�<m-i�jGP��G��4��D
�z��:R�(�.��zwѭ�歬X]^ A���K�S~���l���Ɏq D2#��Rr��6����u�{��a��68�6-�lo�]zPy�<Z����_���[�PP��.�~U����5���8[�f�H����oP/����T��1���H�`���Ƣ�L�	��$�\A}�Z�u�ǏF �C]x�L�yl�A>1bc��,:濓�����s��#�/R�.n{I!+#�@�^�M��6\K6�d��	/~e��*#q	=K���<y.M;K�Y��M�BpS3���p�BW����u�k�jinɮF1�e!�4��0[���bZv��Ĉ`�����hL5|*������ג���5��æIr�ݝ0�YI�gC]e6��ǉVZ}a=В.��BC��ȝ�l'�sP�K?hI������㭿Śb|rݭ�(r�O�v���|����a���}�V9��&���R�����"B���.?��]#5��ܽ�h�2��m#�p��W�飇L��Ž��_�������H@>Rm5��p�T���g+Zm�0����g=�=>��O���F�W�S���>F�F��
�����)֎e��z�)�xT��xy����Y�����Bʦ�����{���j)e�G��0�D��8{C��uf�����	�:k=q��*�D) �V"B�}�W�e����Eh\u:�:�|��(�H�.ryj���<�%\L�M���ӆ����Wn��M^���60r��M�Q:��Rѵ@�f$Ԓ
Y\�F�O}Li���2Dc������Bx~�SO<���s�k<�H������`44iGZհV9G�+y�4ٗ���5�^ƿ�s��X��$��'[9�k_}�=⇰<z����Ƒ#��̊J8a��P8f���Վ��my��|��S���,ci�4� �5�0�$�4����һL*m������A�ך{6��%�{�^�:�"�e������1�O��'�`%��0��;Ic���({k8ݴ���2K�g]�{M�,�M�6��*��s��w�kw+��R����mZ�A'��vr�1x@8-����Fv!:?|�h(T_�(&H#n'�1_]�w��Y��~P������&^�<GŰ����L_�����ݜ~=���k��Ȼ٫^��>��_#�����k�p�&�u�� ��� D*d�,��6�P�E�� �t�p��=�	�D�}1�ƙ�*I/�#��J(S�q��[�S2����IjQ1��9=���mfjU����ZH�G������%��V^ј�Ly�>�ܝ>	ѫO~��6NQ�c..�&j�9�����h��S32~�c���H�Qˆ��_T8�R����t�D��Q`l�\%��Ijɀ�6z�'?���ٓȏ�
�s�F�a��1�D+��`��.����$�iIl";B
=�cjl"�2=��G�$.�1"�'��={�p&�p�&���SO�5���B����5\���9��0�>d�Au�x.:\�U׏<�i����~�\?��zm5��]2.�f�'�]f?l2P��^�9�T����%���&7us^OQ�מ��%�{�n�жc�s�9�l�}��O�"�U-����p=��W�\50~[聳���7߾@�E	��ވS������aM�]3�
B[c�n�\��,����u��F�t��9:;6\�x�������BT���u�|�,)	ۦx�\����+d�4Kj9W�|�5t�9s�ph�%&z�no�� ��hF4B��W��j��(�ZON�3�7?:F�w��&cYޕ��]-�?�;�!Z��c֝�|�m�S�����-&I��g�A2�s}h��z����c���_�+�kv3���4�b�<(˄��r@�I9��#�W��-7���n��(,<s��6�x�v8rκ�#��Ní�57..��������aS�]Zc���4�t���^?G J�P�Bv]1��m.�Ѿ��P;�)�i�=�0�����މ�U�k��F#����A'���r�:KN$!7�]c�6��7��e����t-ZT�K�Z_���f'�Y�J��"]�`��rՀU�gʩ���6M�S��74*0_��D�T+���L(j�Ө��ʯiޣQEEL
C/l�F2��Q�@N�����g�>�R�r�	�k�MY0Pg���ց��y�|:�j�xs����9�dz��<��Us:2��� l����cL.�XGV�(Z&B|��~׮^O7��m�nȊV�7=����8��#���#�-]7�̲���my%,���p�����х%��2�Z�l�E����?#9=`�;"b#4�q[d�̓�%e�``�ճܷ����VX[cT�X(\I�N's-�{�$ʶ�@l�>E�����H�� KBS<Vd��'):��x�.[bۮ>��s���,@�����l�a�=#�pr6@��6��[+i�4�H��"tP�`뫊�\o#�L2j&X��v�R��5c������3��c����y�&�q��ƽ��������'���#fI�M$����ν[u1?`�U#g�Qi38�H�\ϠqV8�)�R/%\�a�_�t3֓���˷9��1(��fv�s�Mf��������4OՍ�|�+Y}h���a��>��H��q��ǆF��̵�@ i���Ƨ�� ]0�p?ѷ'@��3���w�d�$o��w���㘂h�"PQg�6��is���7��'�V�"�o_Xڏ;��=
��2%Cϰ����9z��6望�l���}�x� I�����M�0�5`,:�0����G�h("� �#R��W;���ª89�5��k���F�t�y���k�����v2�%i���c�#�E�Ion���o��F_*N�pސ�$6��GEi4�Pe�I�஀�U̹~���
�"|�"ցPA���F�eT��&��Nh�󭩰����<U1I���k����+G>l��1"�!�Ah��3T������#Ҝo�F)���5�׌|�xί���]��Y��L�)���1��?�vԻ�����?Fi�@��k�E�.dv�5���B`���n\� �� J�Z�ar�ݣ�D>���A��e��J?8w5����'�M����%IED�iinàg87�F�s�Yx!� ����e��\��f��Fᐽb�v��Qb��|t
�5P��o�萩��̅�;g��<d)��K��\
4�6��������t��a��{��`�9;�1�_�9j�
$`gTg��yYOSd'��pڤ<��d�S'���s�ɧ�I���/�skw��6B^z����uѵ�[il����Z�a۲"�&N\�~U2�p�2IN�F%7��D/e��a�2����Z|G��k��N�ߓ��� /�G��mz]ܽ�T�wpO)�l�s�S�%��6�.Q�#'�e�o�KYQ
֞OC�{R�<l��
@D�0��2������6tZ$�"����X!�ա�dTGG���G���i��0���ΜI_��g贇C��{湧�c�!�nl����? 	��1��L���p2n��%���7=�м?ԣ;9 	����pDM��F�a����5 v��أ�8H=�	GF����.�=x(#tTQ��F�H���Z�8Vmh>��`�s���E#�*aia�!��m�cg�^�i2?=^�aD���i6�qX���րE#:�Qz��� $��G':����˷�׿�z�ޤ��{�<���TV�(6��i�5��yT���}ˌ��f�gE�6�KXӃ7�}؃��R�/�g�pŶ��������S+�9�p-sӀ!
� �"���=�=f'��hH�C����rc�B��$��pf)����Y����`�O�v5��������)G�$�xd�IH������:μZ� C�C�}x�Q�mH]o��vz�̉�Eg���;���}i������IJK��s�E��������t����9������wQd��%?),��{�ҙ����}!�RZ4r"�`�d8|jլ��î�ʩQ���e���>ؾ�T3Q.fT�� �`��9s�V?D�,��yP!�pv������]cɚΕ�fT����0����͙R���&g���wlߥ��%�c��^����l�Me��t���6����:���0L�������%�y����AŪ4S�Ϣh�N���W��J ]GN�f��.�������q!�m�[6E;pH��pga��	� �v{��!j�m�*Q�J�����l�:�$����G��%�e�D@B�6V�*��u(���rt��2��P�9�E�s{�����
l���B��׸�<�ΐ2tB��``����Th�OV7��5�#Z祃{'�E�%ŷ��$�h�5�N^��#@��.I����I�q6"�E[lo�z��	�n�Y��H���/s.�t��&i�������~k{�{�EE�,�vg�3�z�å��*bwY�et�@S<��R���hx��
D=�s;L`-�LqP���ٗI'4�U����#�|���Ci��*5��욮ctZ�RpS�u;m���X�h��U<MH`Dæ�lbЈno,K�4�(�!��/>h�牑\[��l���H���'{�����l�2#VPEW(^7�[0ZϾ�*;�"@�
U70�ۢ�ݑ�1fP�i.�����L���eC��)7ZW��x�x��Ml�4���AT�Yo�c��u�}����䕛�E1B�јf4�?�)sL�2}-j��Q�C�}�`�s�;m
8_�����y��ak�K�D�1��r��T�M��.��C������ʤ�8������ہ��A�~�"��q������V:s�%yi��*s�F	U������q��x����=�n���Di;�y�iQ����Y/��y���ʓ���yN+{�̸���P.�G^_�#Í9L�'#����
G�(H�pX��A3-"T��T�F�F£\�Q��>7c INb��#^�gee-MO��L#d����il���Ji4Wxn#*E</��䕄����N�"Z9�"2t+��e�+�>	�Z�yf�&r��@��>��1�lNC
�B��M{HhD%��{I,��3������53���#�5ʸ���r�c�k8_:%�u�6��!�@2?�y<on٦6:��̇���^J4���-׳�sdu���<���e<�la\�H� _�������d�P�O��z4'�����;�j��N��UJՆ���?q4��
�pi5-ݽ͑� �1&z����W�ɞ������}��q�4)T-�[Tc4p����%ZP70���A�:�����{���X�K�ܑ�tˤ���;w6��!m�:S!AD%���#�"vA��"�9�oCi�����D��cGA`���ϴ��VN�O�qe�V;-�Ay<��;���8Ԓ@�C�i�g�׈�T�[�6q���z�F�a����z�dsI*
C]�$��0�f�.�<r���D�ce:�l����w��c��<T�3~W�ij�kier_3��Dd�D���O��	ej��0G5�\#/�0��f� Gu)���X����>4Cx��G�G���ɹIy��������&��0���ڄ��������yY�6��X�j�������\�K?��/FY�5�+��	
������NT#���F����vUY�޹��Ǵ4��8�-�=_Fb�#�	KQj��zp��$*=p`�k�E$�a�����x��m�����-�A�`�<�񭓗4��S5�I� �C���{�^��4]_�����0��6� �MD��D����fD}�s��8�l��ߡ�����?�Cc�uW^C����n��K\ĉ�r�3�'��Ux2�%��o�D�Bڹ�N9sxaKxx<J�p�h�90 Q�OI<rtf�E�D�qޞ]N'���P<>"׼nco��j�e�t6�9P)�8O��*:���lT]hy-�NB(������ ��:�tU�]_>8#��k�nqw�����ge�9��N�;;��D�pҴ�:���EŇ�9�3�v��QG8xVa�Z�j��HS�����a��5H�-.SB@YC���1 X܇�?�!��Gȣc�<'�85�7D��Z׌��P��n�Lgy6���i��ڕk�2�,�ir�����{w���r�����NZ��[Q�"���땕�?�����!@���5 0-x�*�@P��	Q�:|��_�Vk�d˼s�v����0���.�\l�����T�p ��W�;�1��N*"�R� ������cf��O0��Dԡ/��v�11>Q��f�>���Ҡo՚S+k�}���Pe>[�:����E���W���<��M����E�� �R��2����4F�]B�F1�eآ���:�'?V-0A~�K��~�r��cQ��F��<+c�h�,��xz(����z���� �1���gLc
>�٬ȣ>5�3+>7��4l#��"3� Äa)gkWRV��dd��ђ@���� ff� u�B�6�`�E !�����x.5R
UO�/޻�n_}7��W��g?����O��v2}��oQ|/��Fq���k6��!ˍTl�5d��d�l�ns4���j��Lc��U��:�_�>s�ʟ����R7M��!5�;g?�z�sw�<���n/���z���cG�D���������g��:a�:c����,�����w_���qޜ�L9�{�������uS;Z���-�q��N���"<��:>�^��aP��!����2��!}�L`���#ߊ�&�1�w�k���Cc#�},�X8;""���!N���iແkmX4�5�u�N4a�����=�\�=£�I��W��/�V>�(�㒕���l�,�,�ܴ�W-���o�H'FGP�y/��y�Z8g}�U�@T��۔DYjjgƣsm��{���p���M�����1M5��&4�u"v�!�YG�ΐ竓�S��HX��rÒ@�n�U�"�q�B�K���T�7�*�p8�y�%��xpY�W���V"�π��A�h1K$z��7"E׽;Iڃ��g|��M�f���z�x����B�{�W13����uοwO�|���Z���YF^c���ZD����ʜ�t ��ܗ�oB��@�8��6��x��� ߵ�49s�F��&0�>� ��r��t�pO���/�1F�6^��V�S!�`� ���U���^�E`�3��u��UR7nܦ��IFE?���ƑK�鋿NE@�n���
�O�г
��l�Z{7��h}��*��"�1B���������i�=3l�P�h�����٫G��F*c��OE_'B�y-G��{*+RD�����°�$�ap�F�J�]�s��"����%�P�C�Y��J����w�8 cK|��kƤB�4'����PUŧ�'ndc�Bͬ�l"��W�2����0��0鉟�%�P��:��Ɂ]��9/C8<�(5�<�͐��e`���t�&Ց���XJ����ip����o��^yxv-�D8�L2�k�A.P��KG�Q�\��	���;�>��Td���(Q�:��.��&G�1���0w+�L�D�t��Vׁǝ e����t:u�4Uw�ŋ�D/���n��(��W^K�o�u ���<�z�p�vD��.�I�y���������7��T�g��M�WDvP4X"&���4_4!	�g�@\M�խ���H���d_���?|gT�ʡʁ��L{�o�GtS7�E�G$d�^",���<'�N4�tE8�2�Y���nd�=�jF�:WU���%o
F�����-�6��u'T��� �q(�W� ���ذ)�JB����r�lJ�CPӱ��� ���?Fh�h8�.?��;0���Hf%C�c��(��-�c���6���~��q����Q��q��NE�\�X-+S���`��gu��vj4R�����?tD3���U�岭�Q������<��h���e�w�r��b^`�3p6Xۛ��
i�N�΅k�j��2={�b:}��p��JY��	j�-_�;P-�2�7���|$��?�qy^O�@jE6�=�x�̧?Ǆ��N�$[M*,�\á�"�_�߅顙=S�8�߽A�d� EG<�.��K�M���w�T��e�$7�\�y�	�E�e,�;|"��`lh'w-� >����3K���s;P7�p	�w�r���4;a���֜Ħ"���e�v�W��2�7�'з90�ۀ�H	�0�6PZ?���2�yh����'G�t�q�T�OdN��\��pј���HD�gE/f���B�Fj�9�f��Y�u6�D�*���|��<|�s�|_ޚ�<y'B̥j�F��[j4Qh�~�ƌ���W���ε���+��x�6��dss^������W""������|�F����r�<ec��2�r�&hD��Sa�rͮe;Aze�rǝq�ч�{���pŉUF� N-��Dd�c$Ja�5)��'	%6ҕˌ�\%R��O���0lٽL�z񥏧��f�r�N��ݻw��!�Q�}����/>��Iw��vo>r��D������P��W�i�L}��U��G>Ɍ@�h��Y���k�5�ޚ=�(it�'�(nC�l^��������:f#���u Q��%�L����Rh����C�� ;C�ֹ�0���!�n�Q�hp��k[�1����f���qz18��P2_�H�Lsl��$�q�T��t;$Q잰�i��z���16��Q������2()" ���;_�-�����PQ����r��ƻ�f �vߣ)�XP� �)A�/�>�P殐޾�e��s�9F�ꑺ?�kK�jh�U)6ar"��tg�w��*�>��-P	D��Y.�7!����~L��xw����2�)�En
dD�E����M��5�����G�NS�D�����2��!�/�#�lTQ���$|��ie�&�C�_z����c�bބ��0�i6��̮���jS�۱o��UP��n83��4G4�����"���.����	��ҊAU4�a�K�K9�1;<x �qW��'~p������t6H��疧�A��F�
�v	(n�~�>C4��{�h�5�3���O>1�6�0����,6F�v_�m[N3<��]Bl9�Ȇ��w�;Ct�ikhT��1�Y]�hv»Dȯ6���!�����3th��䓶����.CP�[ιE�|��ʨ�e�@����M�#�H��U��aM�e� KY0��[�<`�Z�k>U6N(#�6
6��,�l&��u�G��er����b��_��g��?����_���v��Ѳ���D��Y2�-RX�����r%�\t�:�HL$��m������0�x���k_��2��K/�B6"���]��KW�����/�,$N���|��?������s��HkcT2�+�o�1�h�A�U�ٹ�l��v������Y��A85�U�#Fá�v	#��B8�9��ע�ݵ�@���|�6(�=��a�c($He�^6�ʓ&�
Ľ����W�N�9K*�eR�9z��viM8����,�N�Y��EW8/��т�˳���]�@�۷ɑ����4�\����M�x��-�'��낌���ӏ��4��9�Eo,L�W�}���D��0����
Χ��\���J[�F�{�y8﹄Ní�|uh�f��}),���;�k�qɎR�ו��8�D�[�������cф�M��ӿ	�2���=�0�PD�T+Ɂ�}�7_	o:��ϟ��� ��L�{���Y��3S{�ۙ1��\��Y�
�4�2�=q�i&��K�CJ���GON���Tk�ԏyu���S��[3���f]mw��9����ѧa�ċ ��VV�MiT8��h���􄜪}9tu5��:Ģ3�����Ԓygg�P$�2������t6H��F}ܤ����k�Gwc�O��"0�d-Y�[��O��"��2�@���4�-�9��ذ˛,��y�Uf(3pbַzYO}��J��d��s�ػ*�0�����z#`{LK�臬e����ݦiR� 筍kb؃\����aȵz��:^쇵�ٻ�=����\ë����T������$�қ��ɺ$�lB�L��y=D,�E��=`�
0�P�o���0�:Zk����~����_�b:ql4�i�n��6�Vl���ϳ�m�mY~�W�"�4���#�U6(O�h�X�@�2�����"7Qȶ������'oÌ�9��$=�[o��Ļ�8Y����4��޻7�/����p���V?��v��|ϳj��1�v�4-�9j���r<�%^][��	�<���]p'Jk�P��)�#1��\7�C8�]n�5�|�����G�0�!F.3P��_��)�����X��Ըw9��K���Ɏ�.��9=�����,k�伾�\�C�y���k�F�J�^g�]�Z��c��@%�zzV��0�T�M�<~&��C��!)����ŉ�tn�������[�[B'/F�nai%���u1��ʍ]�<�;ߑGzg��(kW4��k�+k�����~uv�����{��Rr|v�:�=����9����=)�#"j��g]��Ą�]rZ��C������M�F���ˑ> =Y]�?��~p��$A��I.d�p?G�K��ɱ�z�E��p�o��m󩋗.��t��>�&��:��>.18
��ʭ�����tk�;-m���q6��p^�^��?���U�r��??<'��QD�'�5,s�DuFAW6�(X�9<�C6ػR��MY�\�Cg�iY�����V��>�2{�19�i�R<ٻ4sp|��Z�M;+���G��'���7G	T���E��h�ej�/ߴ�f.l75��ҏ��;����t�Qgݔil.Ru�3ી��?TJ�f-��ّ�|�e�ֵIx�φBD����������+?÷*x�K�O��^{���`n��L4}�r��=��a�|cg�L+�s���7�{�aU<X;"u�1A��P�en�&�_�q�@�{_�e��o�GϜrZ�'��2���߇���:���,cN�H|η;�L�u����2����y�
&��'��[�&r]���	�kR�E��#i�p�V�D,{g�#ojd48t,���7碳�5�ѶW�h!fF�|�sDj簬нg:.&#>�,F��	�"��4���I�2J�\mt2��I�C5�6��Z�Q����dα�h&�M��X����S�\�����f+=\>ټ���;����g�_�ŝ�ee���z^wQ{�gu�N;)�g{�K�����r���H?���x�Qq���3!-��Ȋ������T�A�y��q���i���k��GO�����#�P��IH�7��&2#]NH����85�i��`�����D?6�/�k=������?ŋ���={\��ľuUgc��OŦ�t��D�r����&E�6���k�:!��9,":\:���&�lQ�z�>]���>���?����>�� :fvpB\=�;����56['U�5�ҝF�f�����Ϝ�����{w���M'{~s{�4�z`mb�X��D��ٻ�!�{�2W"�o%�m���z&��6��,�>��,;��fC.k�\n��? 	��M�]Cc�#w�]1��'�79����������`s���收1��)���̍��&��f���X��FGzcl�~���=�}�B�R+��w����!�$�{�!�����t�1Wg��a,z�3��?S��:q#+!<��8K�s�����@�R���3R#�؊�� M�+c"[+�l`E[�V=�5���T��F���� �&hD���I�K���u�6�PQyn:FA�˻�B�C�D�1#���LqdO&�hu���O2����+�捛(��8vXm~�FL��1-�<f����{+�:��lUBz?��P�Y��q���覂�=y.�1��ү��6��L(���2�d�0#}��ߌ�Q]��1����_IS�i,���|,o��۟��s�xuh~2�(ݩ$���	_n0cz�p�ZW�t�f6:}���;0���if��P�w�IT��ghN�Y<__�aCVL��c��F3��߸�c$(���^���]�| �Q�����i��K6�����T�����։��= 2�eS���$�t1�0�E8r<�� v'��p��3��!��XG:9�>��Z���Cц�3"c��
���s���ۘ*�x�l�+bd�����L��ؓ|I�t�'�<qB��8�N������s�n���X#�+GS������3b^�Us0��é��J����t͹��ۙ�^��G~>����G+�TF].J��8��V��bg�J����{|��{-�"q�}��{�ôpLf�Fҧ^�T:|`"���I���-�ۋT�D���)e:4���f��H,�~U��Y��"2 y�<�O����Z���]�[Qgz���Nz�:��X�5�������&��p�\{q�Y_��e��,���C�)�����]�����}��m�q�R�5q�>�1�y`]���hM,o��i�v�KP"�JH:����#4r޿o<���!".�쥜i��;W�����~�r��O�gm��K��`�6$	�[ϋ�Р�r�c���<
CtL65�Ad�hc���J!+QרFШk�����5����6`��CDm��ҏ�"��M�Yn�P�PC�j�m��o��A��QJt�&)G"G�hU��%b�,�p��Y�Dğ�ѱ:�����[EL��}�t6�+�92��\�ӷziqy�s�)��
Ghv>xv�3�ȵ�e�����ێq��,�'Tm�lx>��%t��[����9t ���+�����y��O~���ԯ|>�ݻ����{"Ǎ�F�o
����ƫ߂���p����ә��/�QX�'��?�X���t&à_�|9=��Ir��!�����7^M��(������I��W��P	�*Z��o{)1��M\Ѹu���b:4��f�|&Y�)��l��U��@YG����s`6;}<�#B�p��53�Ϟ�wa�ߠ��GN�C��e^m�J��wa緅o-A�p�1��L)��}?d5�*ျ��`ɔ��=���k�uj�,�&�R�:��b D�goL*���d_E~�g��7%�ѫpD�;��09*��!C���mfv�D
��N�4���al~�@��\q����{wn�A0��:m�E�Z� �9��TX���No�:T@��}��p_�#|Z�7�m��de��LTg�GԠC�!�Z�2�zP�&�f'��s���m�'0�q�8���}���Z�m�H�X�y��^��1�N���m?;�9��?ݳ�P�L(з�(�Xq-y�w����0��Ыݴ)��� �)'����U��|�)cOW����8��2cA��䧲��ԘV�!��I�vA^�^�� �{���OA�%X�4)�?0�Ϟ�Cg��k�=[��Y��*OGz�D�s��0�2�F��L?G��3��o~��Z+Ѡarr8��C��8�@�[q	4�&��Y���J�c��ˀ������$W�ln��jt� �$�h�%2i��r><r�U4jS����bw��&6� u�B��WG1Iޱ)���<�>�m
�r�6��k�kr ˊظ���&�`����&kH��*oXfm�� @��2+����Y��C�xB|�-�3���mn>kZI*��S����];9�0X� ���rL:c�D�#�[y��U<:�q^9Z��q����ϾU���Vz3�:�����0n/<�4p$9��A�/�6���4�$�ur�+���(�S�O��|�s�}HE�%���Nљ����~?Z���N{��SG�q�'�Z�;W���K���0�l��&��ߌ)V���8���o���H\����܁JI�P�x��L:s� }��F�߫�&]���a�v�k�_aJ��Y�_��K�yr�v���u{?MEΤ�Qg�w�{@��K���l�B"d
�k��/��Ȥ6��8ՃY^9v�f�/��lKk�0O��X���<R�=*�����Ǡ�3O��9R뼯S��Z��{���=��$��lr�<Q�E��;�p��M�����c���2���7�E���4���>,�ÈY{�kū^.yz��B��l���^z�����
.3q6�KQ�k�ܸ�O��T�ߓ��>���@A��F��+?�?z����S�D�b���CSp�@u2�C��o$�.m�Jdx#Cަ l%\��q����g�����O���p|T؆~S�h��q�
t(;k>���A��d7���"&[h�����p|NJ�p�C���Q����v<���.H�}���A�� �"4��>�2��$�IY�8��+���� ��$��?�<d�}(�i�n.�)t,��45�(�"�F�KݩZ���^D�P����؎,ʦ��5j,~��"���%Ym�F�vt
�3:y���vvw#s6hg8�Nm��WU��Ҍ�A] i�ƏA0��e�Npo���L��L�"����
�L�k�����AP�",��D�]X�hacx��NBVO��a(Ҽ��R֥�|D�����a���_ߧ���)�M���#}0D���،�H#>��i�� ��A�
�(���5
��Un(���s�թ]h"����W��M�<���*�����L�Pɏm�$��q"�P��nnC�i��#L��3��;�Ӯw��>h�׾�=zso ����󏦓����cy�����g���b�H�	s+KK��|�f/"���Z��� i?�;�u0�#�r��W��g�{6=��@���}#�\�s?vx?���� ��6M>�H�MO��{�ݨ��_�?�������/xe��ԘQ����p�z���`׆�l0��Y���R�~+�'�����m���E?!��`��,�Zc񆬄s���C�p���h��u�|Y�{�jq�ϻk���������GX�t.�b_��N�cD�sG��ßX_�5�#��8`�m��y?��FV���g!�7P����'"�
�p��3��*t����NA6��{���do!z*DE���ڬ+&)
=�&�fY�����N8s�Zg�9L���@T��@�X��<u�C�����y�=W��q��94������Wq��d���%�T�x�ڝ��#��B@)���@��0��I	��s��� @<R�`�S+ {p�Y�SZz�n�̫�T&�6���i�;��6��,�#�S�"�-��9Ň*Bg�t�q~����(w��B���Sȶ�̃�@�كD�ܓ��ai��Ju��R��*�@);[y��l�hroV�yb�~���i�~���;�����IT6�aQjt���p�V�"���bx�z���*#�MSe�X��f��˦��2Y�1}���],��� 5�[{�
Kj}�پ�l�N�p���(�ql_iu]��\�΂�D p��'��gTFA$s�n��+�ȳ�v�!��%�5���W���FF��[�*�_����N��d{�L��Z�P���!!eeyTϗ�m��}�J�v�oM`&��(.��W��{��Eo�6{�e�Ca}�Ԟ�t���t����vz�߇��wd%t�Q��o�}�$�� !a|ǐ�� i�`�m�Fi�O�����\�.��;���o�St|���(�Y��I���`��"=�'=M[کt�� ���hR;<`�܈>ܤ��?{�aK��Q�{>G�x��QYb��̞�J�����H^�|�9�p�ǿ���Ty��A`�A��џ��'�3��ȸVｋ�{�b���q��/��1�'[�p����+ rƳ���ka�#*��8h�v��1x>O̟�$���;?�?�Э���ڳ�K7漚=VnD�<�u�p�@؋b'kP���_�l���N�<�`H�:Ƭ�d2�t��edM�6��и��&c�DT�a�M��+ȸ����<�,��'ݻ���@����iehYÕ}��0�#�u�0�Fy�~:b�0�{Z�/�
�Kmܷ����-]mP��Ŭ�v]E�
?Y��bTW���:7:�2�Ȉ'F�ʠ ����Ed�z��h�@⦑���ׅ�
n���Y������F�F&"���A{ L�0ǲA+�#����	�I������l>��-�Q�ލB����z��P�A�����������.�b��0�@mc�3�-��F]M#0\�y���U���ı�t�:}��! ��?�n�74'HT9{��J���MI{��r���è2�'V*��yؖ�mn,��$��ڦ��D�3�14�Qà�����
ύ =�����#J�hݺжd4Ks`#c�������U(�g����^%,�%�ĭay^@��d�K�3���/�Ґ�R���<:P�:����az��U�9�o_yI�S�E[�BۍzY��k�s���pUA����5��Q\���M�=Ӥ"��[�d�hY:$2��ޤ��n�=���qj#�O۝.�OP�+3���|� �|���xX�Tl"� T�M��2�m�ק�YYZ�8><��.��FI4��K?�Ŵ�z��7K�9�f�&0���w����:��:p.�Ƀ7@	��A������.�� Ֆ�q�w�Thݟ��3��9r�X�ε�i�i:oi�HX2�萐�3�g<�lbd�7�����XVs@��F��.{��Y"as���b�U�W�W�OAZ������5t]v����,�L�|u���gr����8����p�>q}{�#�C�Ĭ:�Y��.,͑�ѐ��aw����9ɭr��"h3�Bגh��x�و�o�uep��67Wu�kF幚!� �!;��8�p�u��^	�<"|��93�!S>�?�1z��
�6�n|����[ A����:e��?�� ��P����kbf3����~by��L��nz�����HW�K#za�@.4��o�uw��]�/�reN�z#��ѾF��z��H������{=�9��-���!Cfɽ�F3�2�n����K�%؆#B������
3h���1Ɔh� �Q&.��_�AgJ������[;��l�L����H��z��b�W[�v��"�i��o��7���{�`'��cG`$o�ӏ�:3Z����E|u�'}�{�h�@4)�4c�a�l��B�@bð�O�ׂ����U����	�L��RU�X҃��:#!s˧��*}�."9qg�)�~�J8	#�*j�e��ǎr ��]�_�#�%��������oGF���ɪ�)�b4��(����jF��䒤�$���i�x�|�ǳ�@&�6���^fԢ c4�iёМ���ܣ����x"�;���w��=LO?�D�Y��V�ַ�G�c8��t�*���{�v��I��p�.Uw��%��{�4��q۠]h�Wei���~�f+��F�Ʌ߾7����8x��>~:�o2Z�֯2�㷿�C8��z�J�}���6h�{c1Dk�:��L�:7zV ���xf�B�]:KDB��KD�A��ܹ� ��]��n`�/�܇.08f��?i��=w!���!����?��QO�"<ʄ�/|�Ӯ `��i�|��<��c�,���w.�7'�=�]C�a��t"!��@'Ѕ�m��c�/�oF���a�"ES��X�F|� �[��p'��������Wk9���a%w��S����v�NI�����=&�]�p��q=���'(C�q6��~;��Dݠ��:N��a�����u�a\�_εߛ�S89w0����-G�}�w`���ՙt]C���-|-�/��:�׍6E�D�L4pny��o�r	�:�NST�A�����H�]&8����gi�t�5�7-�W"�蟜	�r�D�D�b/���Yg�z��U4����U��Pz���u�H@��Zv<"?����E�p�E,�Y<�u(�ևS��R�Mw�+!�	�_����[��ro*:F[[��ܐ*ΩVԃ��2�(�����#�p�U�����?��KQ�:w�,��h:vd����z.�����p|b�N�m�k������ŵt�v3ݞw�'��
1�x�6f�[��t��jqv�I"��� ǵ#l.�\wn����&������(':�<e��=Bl��Xv�<Wgoս*^�\�ZMC��
'��n����8�0�UC�N���6eG��@���%k�&�5c�9UZYA���x�+�ʫ�%��r^�a������6�Չ�܌6�0���y�w\T�11���?�����NG]��O?�^z�t�|�v,.��?�����D[�ҋ�?��;{�'�>!�w��q:�Nw�F�ۿ�?ŀ����C'�.d�y�][�"����0��?=�R�09�3�.��}�t���4��Yy"���� z���-������\��XZhn/p�}�{��$Ұyɱc����x$���^Т���D��S���]8�~p1��Ǳ�nݙ֧���������i�=�y��U&�-��}��P�|�4�i�ɹv�l-M$bB	���O3&lU���Up�En%�M�$���ôLV�n9��Ʈ�3�����F�ZaP:uВ�������\�w�F�:�fFJ��v�15C��ԑH�}p�F8k5��6?vvfo�!3�Ն;`^>�Y�A�זIk�����5�{\���:|�0��~��Aw��{�@$tIuݺ����aC��R�$�^�)B5Gr���1�3�s�D�r�&&��K�p\���w�)��vA�Vl��J����L�	GOlRn���hiIe-�5\�����wx������N���%ջ�$��L��_$g\/YSŏr
��C��.%��|��@"E�gb���W���U�Om�	8,V3�07�Rb������2��f{x��;#8�V�1�yǘ����1���l�������(]��uX�F���PZܐ���������nݣԫmH�gK�-��<WV�y��l�a��#h�S��ˑ�Ng��Cx��|������9��r ��ψZ�Q�-�'�.s}f,lK]�n���*��Mf-��I�B��Zd=���������/�,�GVN��*+��̤��=tx�묈|�oGO�
��$�Y.g-�O��c�c�B鴄��X*M��lb��A� bt�0�w2��z#?z,r�����ӝ[7ҋ�=��"ߋ����-����W�h������O��D���>BW�u�rHJ��p����W��jL_3��2վ��_��U��%���4E���%�t:)!���#F�j�̢�eV����`�׼8܎��uo+��W~/�w�c.��GOГz��=��J?Bx"a@����1��;����?�"���߭��t�&��t��.��$�i��t�@&L�Ds�Y�f#V=B�C�x�DǱ��;
���}�U���Q�r�*�F�� V[�b��*���3h�+��oTgh���1H��Y���eHf�|�޽;��7���3U�׮�� ��A�(�1D�"��1��=H���q�c��G�uF���8��i)sǞY��Ξ'(�;������G&v~h���y0~@=�g;L�
G�ja�m̺0��w�s�ߛ���,�
H����ӧ`��`��.=�#���e�~�x;-o����!����Mp.2��9׏NN<�I^S�f=�s�BNdl����JF=*g2����#=�w� ���49oT/z#��E1x�T\|&�r��nҒd<��b�����ԛ;c�����9��(#ٻG?9�ç��ZIo]&g[3�:��܏��Kts/]��L�r=ͭ�E<�-r������<{��wQ��˟��s��V��2���g<jy�.�朢	K�7��7Dd�r��_1�H���{������N��6ca��=�P���G�֫u�&.�rbSDUYɆ�ז�]�����\^�P����|c�ge��ZF<�S��C �\ͣ�����x�U�2clC�B����su䄉�Ǧ���(�A��w`:}��X��W_al�Uƕ>�N=�(���LG��Д��Ё�fT+ghA���O`�oG��g�|"��|�;���$���215��k4��|�m�{�=�Tc��Q�*9��qmsvuIH�s4��.uP��)��ӽ2�;�;���!�Ћ��(�e?��_��m]N�<'Ym��w�ʍ��k�s��w��3��~�!�1��{dO�z=OP��eX�0�(IE���ɐ�=F0v,S�1�&�ڽ_�{��B��:�r�����A<����Z���u�n���������:��D�NZ���A�;�'OF�!��X��k�15��"��ӧc�mo����jz��+�7���vY�2�}C8�:Y� :Q͜��p��b���\RVE�q�dG<�@�V��E`lܓ}�Q	ע��J'�c�uz��{O�}���@ڂ�"o�뉮{8F��8i;����A�γ��d�-�8��q�M�&�#���YƧ�A��nI5Ys�`��&��<��������{�-�MF��k�ㄇ�����YEϡ2>�O�'��Z����\)>g����?�Az|`ԣ�:3Ғҗ�@�؇�L�c����>�m���������C����0�b������CE�2u�M��`Eұh�n��Ǿ�ɦ1]�FD/b�@$�bstl�wK��Rm���Unz�SE�|�����z�18�����aZ�a7�}72<�܉.��P&����KS���W���;!��/�����99�*��Ȟvg����=��
���k~8>_p�e��>��v������Q��<6 �5�iD$��.F�Un4�N?rA�41���	m����r_x��K��s�1��ߩ�Hw:q�D��'_�П������(�1�3zy�շҟ|�;��Q`1%M��%?7�\Ow6nS�l�=��k]#"'�߻����@�*���W(��E2�\*�D߂p����<9�=�������;2E����O�yL79r����z�c�Pi��q��8����X?7GE�:�~�.e< ȋ�B��AO����e��j6(y�P�����S;rԕs��YH[G���0,������d磏���g���r3>�Z^XqjJ��w�]�r�UI�rb�TFGgϩgN�k��RF�.���:jM"��1}W����4�F���n��j}�pƵv}v��$�lУ�Se�;<��;0��r�[��p��6�;\Qy�X|ǱN7Ea��~�J�����UxX�c���6�����Q��2�\�._��M���K�}�\�U��j8�̛���T�s��^��*C����x�����3*7�/G�!��daf'�k�<�̉�qs�����]XX���0���c	�#��O�Z���`л0��]l�c"td`��z��S�?�)R�X�5f�I���9T�M���a-��N�nE�9JeQP�m8��2;Dh�����=�5pvd,iՈ����Z�����z�����؅����U6|��,���Goǹj)W['+��wB1�"?�sN=��{$�Ă���+w�D��9-s�:��#�9 aeӁO3K�s����U]�����|^�;9��>x� V�e��T�*�0����ʴI����e�ixQ���w�yV�Tٻ����"<�T�A�Wh�ڇ����^���>����Z�I����7ކ47�����}�#v6��r���4�y����W^���PA��O�	 E��5���j��MJ� �շ�`�9l���E��;V���tTp����:�p��T�_��g(�;LT����ۯ��:k�DGP�An|��EW@�VF�ȉNd=}�{����ch�Ҍ�� fņA_� �ʶA���	q܀�JU�sސ=0��p�S�y����S�r��j=U�6�!:���笸3��y�Y��1���mB����3���Ig1b5�μ��b9�ߧ�ߊ	T̌BR<	�!&��0^�}Q����:�����N�� �g��'L�/��N�;��W@1��,�����=�l�G�����`�ee�w�6��3� a�)�B�K�6*�s��7b`�|p�\�ѱ�#8g%]�v�~�4r�D:���c�+kd�VŐ@���Xi"J�>;o���k%�]�*���S��*_x�GF�᧕G�}��W��B��AB�9ɜ�xs|�����s1_�ȡ�8+��vA� zF�*�K7��U�����{�܄������C��y�����Fz؍�#�L�Ƚ�BpI�ǅb��#*��v4"�ګ��,�Ie�����bA��9B5���$6��Lk@�Q��k.������jE	7R�,�݀�9'TO��ig:L�����@z�-�N�f�=��lO�#R)�8��\ܒ�Ā�ܐ���{�9�������&׸h]r�\����]U?e[{f �Y��ʌ�DB�֝�ˮ^Y��>[������85���9d>C)���n\e���7�Ï *�^����O�lS�x.���+� �gYK����(��i�Z��p��\'im|Da�*����fA�~n4(��1���@?�#�����*��೪%��!D�f��W-}�� ��H���3L������R�o����Tjo�%��Q����*��cS�H5i�@k�m���s�' b6Q|"2�:'8>��^wJ� �+��1g���c?i���$�h
aJR�m�o�IÔumg]e�e���R)��?4�Y!w:�uT�e��]�Iվ	�?V�Qn�~}�{͙+݊ ��~�\!�<�z�˙'�Nئ����<�T���^����ٍ9���7ixt;"^�"�̺W�UT-�56y�_*yT�����bLj<���3�7_UE�_9�g����S�q=љ�����`l��Rtb��w��1ཬ9�� s��4��_����Ѿ�N�

�E����r �-�p��,�2Б�"������f�iaD���k���2�A�
LG��"x��sّa�ǀYt^3"�<w��m���ܼ�F�g1H����\�^ӊl�%��^��'E��w`�D�y��D?D�����6�+��<���(6���(E�Xfh̝�4�"Q�e�I��zn�|7� ���š�7W����G�0:��%Nؕ��.C��
jx���Z~�JFff.��j������#����^�$:{R�$�p;-c��$+լ[��+�"_V�0�1ؘΛ��7Pp}||�#���UJ�~�Ыt�v��e��0��&N��]�(��%\��X[[F�[�x/g��OP�.������Y!𐚊D%iŅqa��LO�>�����s9qЌ������Q�(y��~�Ԗ�#/��y�0�E�-��_���.o:*�]deXUu�Mt�˽�EO�:�'�{
�����?�ĉD�����W���w���f��=F{U; jX$�<j	���ko�|��-"�z:��.�=��=�}��W��^c}�ZE�8���h��z�o�!�!&�� d�ē�=���^!�aJ}����%r��0��z�Z�.2�n!�?��O3qk��R����8߽���|�|����a�4@�4���!:ު��Ó�ԇU��L��Z��:��H'���X9�<�NGC���u΃8*vb���"
s��SM?U%�UE�L܇<N�P�mR��C��'_�x:)ν:q�����\���2w�u��W�Z��e��c�����O=`��r�'l���gL�䎇:9��R�A�c�s��Ge�#�w�Ȗ��&a��K�u����z�)�².?a����8��L� ��6�m�{��{���D4���mrYo�/$�Z���MR�C���dnBv���������2��!(�j�N���e���Ι!O�����
I�`���)�84l~P�T��f�	U�,�j0@�1�|�~x}�hܻ{Z4br'|ɇ|�M����u��7/_e|�Q��Kn>IsI��1z�x�uGO������$6�T]p*L��c�.�M�RjU����xWRq06c�қ_�1��9�pO�$&��ػ�m��Oe���>[�0Φ|r��f����K��zoTrT�&~�y;ޯM2r�'�gE���l�_D]�kV�U�@x��<d'ō��������~"�)*
��9��g��]kN�����T�0m���5�}�א{�g��<X���'��C��o��oR~8��i���<s�Ӕ�����iﾙh���_�ٴ��1(f��@|z(���ϒ�勃WW��s��5�����K#=rpo�s�\�����rg��6D5[hv�s�v+�t�γа4�g�<R*��E.���}������@9�c9G�O}�3��'ǁ��0b��̠:0�o��?������1z�?��#UyR���;\Wo�؋�F�L����~��ڃ�DZ�t����[x��Q"�����}Ϝ�xl��P�9����עL�E针��hB>qo�>��������Jp/�1���b}���(h��J?�Qw�屫���uHe:!F�ƛ��N󘈘��N���\f	��1E#��{��S!�e�)c-�2ט���or���0n�Ͼ�zD�y��g�d�v�GE����1�E]�a ��>2r�7��H9�;)�%����v._FF*�M����Rb��i�=��=�#�>�v���V5�IY���W��N���\"��$��9�t�%z}T�x�����M�}��i��+"W�A�m` c3F��t��n
nQD�o=�7X~o��`�	���d=S!�ٽ���2�to��R�5J=oA�=Js�Q��V��w�R�I���!����d+<��L�z �A'���\ۜj��vix�)��n^+o0�R"¦q��Q��n&��m�����=�~�?�<6�C���v�7�=L��##Мc�SU��U�gD���=K/���22��5��5>�V sw�S�;+�e_i!v��ߕv��.���9O�6�hW�b�U�|�{*�:o@�5;��d:�';���4�p���_E,�/vf'2�0��:Vt�2�y"j� z�1E��^��D5�K:�܆�r��vb��;�g4:~yO�x��pxV!�&/nt�3܈�0=�3DgG��ƭk4~���a�v�/�����
t'�	��NPw��ϿH�j:���\(���at8�۾J_�e��u�Ɩ�Q���7�z4r��>��:y�<C~'��Q�H������1��ҥ��������ν�V�'Ϥ=�G]���bf�,���xz��gXd	1rO�\��M�q�f2�~,}�ܫ�3���~�MӐ�"�-���ٗ�L�	��L��A<ξ�A�x}���{�[��׿�o�ЧH��M%�7�u �j�(�[LU˨���Ԙ+ha_ｈ�#�Τ�\�.�$�aV�ѧ��,s�����Q�[�*�ؽ�t9'��X3���Ǟ8��x�D6��äh9�C�҅�OV���"��f4����� ǏReџΞ=O�M�Sj~�j�^��;Nx�q:��p��\ّIpվ���2�ɹ�<��=�EO�)�㾈���\�y˾`m	)w����8c�{pY�8�ΤXY��w�����G�3u�	(�&�<w�6�����i/e�Q�z�Ug���8�a�=�̯��Cu䫏uQy���_�Z��#b{[��z˺!沮O.�Xx��0��>��M7��g���O�+��!��UĔ����v��£���Ҍ�F̬�<V���"q� ��� K'XN�&�ue�\0F�14��25�2��W�8�
���ƊP6BL}�L��S�8CfC?�z���R��F��Ӽ�s���vʛ'� *���Zc�:G�Y��66���q�\�c<sj^�d�^Lw��Oލ�:Ƽ��$d��#�/�떍�4��)=OٵC�5'+��Ӷ�F��(���!���^_��J�J�a�g;E�i�s�������t\3M1��=~�P�E�_�cXI�t���۠��.�@��]"�4`�{(9s�N�����0�ֆ��]�z>���l5m,�M��ۿ�W�2��l����C]�a�F���{��p/�9�#N��S��ؓ}��XB��sr���>_x��������9i殹x���0���|��t������a�k�+i?��Ǟ|T
�HS�����t��Y:�O߄D8	j2̐�	j�u<��>7V���ܽ��9�pEkQﵭEM�X�o�ܞ藞SP�|�<�F�[5�lU�fX�hm�i��a˫4���u�i�KT���h�i�{�aF���Y���pax�(i�ҿ��c2�u;�T�"�#�FbV�
|�\�!$t��ѕ��4��Ng�r̟��'�k�x����-��������Ty�d9o��\G�0��5���ӂ��$�'��@0��}{銈,u�61b6��V�L��ƷM'9;��]��o7���Q����"��R��4"�7��C����\3�BʽXom;?�)�6%���z.�HTܛ�;��<T�B�K�Lv�z&�z Q��^�ϋnMG_����)����T~OF�2A�~��3�� �[b�i�]���q�7�х{�� �n��*%W-���Cd�wz׷j̀{5Sz�n"���hّKғy^K�r����܌ja廜�Ю�
N�Dr����gr��e���4Z��!��&6Xz���������+��+\�L��(8|��l�c�g딬��.e۫FN<�ad��U^mؼ�H\g�#�!d���|�I��"w�W�һ`����1ר9)��~�^��4p��޷o߉}�zn��5�,7����N��L�%*3��ԟ�o�FqF���T�]�M�՛W�+�~�aY��`������n�Ay�մ��,+�q|�ľ��g�A��8���5R�ְ3�3�R8�C���?�v R�c����F׷��qbRTUde���i`t��O�D�^K�����rm���̜t�A��W����?�����E���0��j|���v��W��t�#Np{.=KıB��2��ƨG�vȈ9�l��aZcMi��0���V�^��� ���a^��w�UGe���xUד�x�f.��\���^��N����bY��A�V��%v:z�No#�h�:��$#j�W*�ƿ|]΅ǎnp�1G�9��aSO�@�b� �G����h{;<2��6��=06�D�;�\%ne�F	��H��d$s�;w���1�<cT/]�2�^OҨ��k�+l����Q�X��`������V��A;u�"ts�}C3�I�K����y�Fs�Uk0w��с�B�;@��M�_�Be���M��} .�v��6�ݻ�:����،�>���9���c��*�nm�!)I����ʂ��d��y:9��r:ݔ��oP�Fi�h���_��p�\[�@��^��}d�'�x�5k�u>TU�Ik;��\�:p�|?��)ҡ�!��m��>���C�?:v��3�@Vԕ��%w���aγ�OF?��b:Pp7�p�W0�9_Vh,3^,ܜ�	D�Y�*����VT�BCAt��m,�]lP�U�����2�ݏ�>����q���UN/�E�m��r9��(�.�������o�`^T�~��mY�v�y���-s�*Ԫ����ݎ[ű�$6�p�"�-�f��"��%��g������#�9��:o�v:56=��ݲ�Py��F=�nA�@�lA�o^����׾G�mO4��x�YF�j#.�֏S�"W�L�F����"��)Ubf���d��"����`�����~"��ܩ��[o�{���W������G��Q�1	AU��s5񛪈ҿ��s�YAi���Z�����J����~��`��4|+��o�)��'q���L�1�w��)��u�Ht3�U������1�O�!:����i��;��`y��ōk���Z�=��9�����VV��=�XN��z���(STũ��r��N.!��*gV�1T'��i�Nw4��gGT�-:�5���,5t�i2	M��r&y�-#�����|�e�a�������g��m�o߾��x� x|���x%��x<G��i�$� ���2��*������'�y��tz���A�He@��Y�Zx���2F��wD�Az$�M���B�Rk�0�+�8�D��ip��	s�7q�MMeҠ����u��Ȉ��#Jg����qvGA~N�<IJ��{��Co����bOLl�y�.�hG�,�auD����࿄!6�s�s�N�0|>��R��5�x���1P��`91�j�����Z/Q����B)�>��1�zf�ğL��] Z�Xu ����0ʬ��A}<4����=ֶ,�d+O1"L�ܬ|\���'y��^�s^u<Q�Jt<�Ji�W��>��Ex����A;�r�&ǥ����v�r�F�� 	�!:�5�@#&��aFw�~q���+%kE�<Ɨ�AI�	;������r#�|����!������h��Fj���yɡ�Sn��|�}�g!��2��_�x)ݡ�:9m�k�C��n�i�e�l��^~�&�P��dUO���Ї|�(��.ڵAI�6��'_�z�����)�sD������ݝg��
�|�ȟcحrDaF�J��z���۩���tg~�{���;�+�d5������Ì����#�NyM8V�֨��/���P�\�����t�����@�0��o}�[1(�5o�O}�S�I:�E-2�W�thd�(b���4����=���֭t��Cm{�6���;�������R�iQ���fz��7 %����G�o�
܄W�5��v�����M	�~��)���ʱ����Ga�-�]ű�A�f��鞸�9����p`b��:�EB�Q&���/׍{�cu��e���e� �?oC����[U ��g@9 ����q�y���C����h�kt�T�w�Q˽"J���8u�T����v��`Ȼ�5(Ά�ꢪl�	�#b�,rR��O%�Ÿ�j��%q�������_��ݼy�gv�:�"���>�qtC����-Ċ�X�������@�,�?p(ƞ�q�LL�q����=��R��{8��_#��>����=�!��{4��%���<�.G���r��+~:v9&6O�d�T�5���>�1p��Z��qo��Y�(C���p�n߼�=s�* +�q��Sʺ�A����G4���} �����zsd{�5��޷�|�V�aHd�g8.TQ�����\�QAE�w8��#z�Е
�u@Lya����.`��3ѝq�전>B��\��H61��t~�R��s��;���5�l�ةw�܇!H��(d�f�s�Jиg�2	$"P��弝LV_������%�F8G1Fy���۾��,�~�4�H��6�O,W"���(���Q�K!j^U��ёp�o G���K����(��/s�{����U �{�΍��P�f�,�I=���Ŷ������u��u�r��j�NR(��A����qZ O�&�/~��4��>gڿ��;��D~)�о���G6>2�u�$����r+�[4��mm�
������'N�Z�D�k_��{�6���F^�����*���A����~�k�FIΥ;(y��z�V7�D�<}8������H��_���,�sm]0�q�������O}2}��[����c�ƹ��&�K��3�r�bz��m=��\<s����sl3�r��ͮJ��k����7��#`6�y���T��8P}B�U���a���ltɑ0w�~׶�QD�D��i�+��:�F6�=���N���s|��4��=~�h|pb��2\��;9p���H+ؒx��Gi�j/������e�IwVh,1��W^#�s�>O�� &�  @߿z�%�r�E�<cxWWX���:�4jqo��c��Q<�W4�1�䵍��Q������V _�!_���L�o��0��pY�Ni4�721�1���>;{�lZ�w;}�/��g~�i2�3��@<ۅ῞��!	�[�����:�a�ÜD_W�J�u�Gu��J?�U�&F4�S����Bh��D��^a��>��Y�RNG)�,M]B�����Ξ+�h�O�9U�;�Ý���~P���t�0��z1LyZW^�y��R��Zbmi�ss�
�*��X`�T3��s��s���y[�����To�����a�6� `��h�R͜��ߕqvJ��p_�g���q��Q�^q�$�Ԇ���mw7cH�4c�8��k�P�tB�Bn������b��%�H��R�9J��4�*��(���F�����Wc.Ԯ"�3�N��FG���*�W��U�v3�0m҆U��Qo�?�s!�EJR��]��)5R66�X���ܺP���T��wL�����'�Dc�e��m]� ��l��wD#�Ӈ2�(�-#�1��.�O��L�obh���{<=�{�y�_��o�*���P�Y���0τ��S���Q���K�^cr�ݯd/ۀG�A�f��L�r2R�V����9��ˠ᡼!%:d���b�{h�W��e�*�>������˫�1t�ֽ�t����?�7=��)��D�sN�Wg��O|�}���R&��B�m��a�<k���Z���:<N��9e�?�����/�wY�N�N��d_���[��7r5�y�㸹ǁ�u�c	��6`��TG�q�%܃N^G��#���
���rg�B�|�.�������KW��7�#�� ���k���v����9u���7�*�q������ud����s�3�k8k�������X~������$�p��?�K���͕�쉼u�χ�/���sI���\(�s�8-����8��^p]�~(�]G`��;�1r���Pj���Y!�S�|�Bb����Wz@�~V>Sv�ׅ�="�7Dֽվ��f�����W�B�ބ�rCx`0n=�J��=T���8	�;oE:Y!=���Ơs�v[u!��nN�d{�s���UD�`L�A� h��1�ܼF�z���_8x*��Sv�l��u6]�����X�kHr��:�4���d�p386`�L��	X�����ߟ�B:�Tb�x:�6ŀq����R���t�#sڈ��`��W��f��@�疙9��EW]E�ѣ>�Ϡ(�G�d/��.@�$4{�ˆ^ �Q�h���c�����yB���-���]�m�n�7ڐql�5�FLAH2B�����;i�!�^��D�^�~.a��M��oI���F�J�KKx��a"�IF�.m8"���瘔5Չƛ�+igdb�i|��E����N�,�:�=ޭ���T��}��f����(��R�v��8"k˞j[s����0"�hʽ|��q����v�zI���_}����uF���ޤLO��#����Z�^���ι���}7R��ƶx�A
�,#TW�G��n`�q�~��E΅��{��a6s$�ݢ�o���ƽ��^h"̽���1V=����Mk ��W�/П�繺CC�w����- Q��0$��L����@f��2G��GNEU�0��~�m��o}땪�RU������]H���Q�Đ��K���L�N�n��R�E����;T[�u�%�����Z�b歍�={���7���J�"tZM�,c��B��w� )�)��H佽�؛샚�hN�!u;˶�8��:D��$龱W�U$"��Ȝ�N�!t�"r0��c*B�hG��Bg��3�r-l�ZR+��mЦ�_�~:��I�H{�y��.`'���;���[�hdu��ߟS#��*8���s��\��0��������&;��p ��|�Y��誟*m�P M��|ti�5��Q���z��0H.}�~J�6�����ͭ�16!61{�>bL%"�Xe.*����Z�MP�D�l)�c�C;w�#�[�6�ϡLʙ��t��F+����&����b�Z�eF�1N3�����N���'�/_J��*j#��P�vF�F�Swʦ6'��ly��1Ց�$�P�Q�A���	D'�$a�rI�Fh%21�l�YX�C����U�[o.t��{d�˼�4�1�nr�d!	J���Їu�4c�s,��m)�{��t��T�'�wӣ'�{���/<e7�w6]���g?�I�?�z'����&��� �>r0����+o�M\	��nh-��/�җ���@�z��(�:�b4E�a,<,�1�]�k@h4�7�K��VwHq�KU|*������_���@�1������|��my.�X��'N�"�M�Xk$]8w�c�� ��v��(1�m��SGN2`7Xn�]J��o�Q�j�s����15��8�z2%��,�}���t#Ƞ��>������r�i�k��� H�����_������d��&�[L����!+Z��,p#kj�W��_�W�b��K/dh�{���o���?�/"���Fp_f?�Q�(#l1}�3R���7߁}~!]ۼ{�9�O����K���^���������	62�.Bg�"~ s�k�*�o���y�����1.��"���7�*�f;3�]�̙�w��x}F�����}�����{�W�/Goź�=�@���[}�S�;oaۙ��zq��H)�][���bE����r�}���>�_���;�O�O�g/�eV���mP��`F�L�I���r�W�{':��[Q���C��S����e�<� �Fu��-��:D����>����οh]�K��*����{�4J�U0R0"#��A�F'Ӟ�T􊸄�������t6a�&����F3s/�IwX���4lq��ш��N��J7W�?Ls��\T�N�yf(��+c6�cpUFl&�f#P�������-ꞷP�}���N�G�,��+*RHo� �|d�#��pݢfya�u6�i�U�g�"-qst�g��7�-�w4d�Ǿ%oY���������㘟q��(d/�9?�۷`�Z[-\xY���cR�
�s��(�Y��;�k��F��Q��J���{�3z׸�6��Ds�(�1"뀾Q>W�m�t����%�3ju�f)F���[0��hr�\�w�|�hMp.��ޚ��i�r��ݺql.=v��������=��Y�S%Z���L�j�b��sS�,׌���H(uv��U-:\M����D�C(�}����}�u3�޿L� �e�Gg���~`Rr�������T,Ҥ����sms9zD�`^[V �J���A�K��k��;>�D�4�	'�{0 )O�Ns5��7"�?�ǁ����8�g��뷙5�à�aCU�&�ڒÉ�	�O ���#���w���������N���sW��>s�t�C�C����~�Y7�����}M{2��n3,giy;���p�W)a޿E��.�>��6i��6dɨ��Xc��_A��$E-�k�r8�h	x� 2C�*���"`�k#Ĝ�nw�t�-�M���+Y�nv�<���]�Y{F�~�id��������0�w�6����kئlԡ4�� ��O��i��8�i��7�x�4��4J��C��`�qFYU	�|N�T���42�ѹ*2�x~.;"�b���&4�C���c�Q����N��o�L.�X<>��!��^��cjѲz9n<�Q�Cc��J�t����7�n���$���m������hT��H*o2�d	:�����qF	�1�10/�XX������S;0u�BnӃ
��^�*���DL�I<6��nu��jy67��;d���d�8���sΞ��N{%L�n�sf��,�$b8=r_y�Z�[��A�lAL3����;G���Q�؅c��ߛ�]cn�a>3V���!�k`��ڐQ���(�c��Z�񝷧'�ϫ��v�1$��K^�ƍ����(x�M�%ʙ�B��IG0����K�>�,p�X�G�<�V(͙�&ơ"�H ���"���ppT�ܛ��B^�I�h"��0���^Φ;�<Ɍr�A�qm�R��֮�(>�;�Ǡ���+�џ��1�ͨq��>��t�Ң���:z�<�8�����*�D7(Q#eC��Q�QyW�t|ns�4��q��>x -��$-ɗ$�__�&�2nL��������ԏ37�3H��;LΛk��ܐ���a�9���Dz��' ꑣ�fr�鐺�K�	�a��l����Gy2���O��Y�|��)�D��Zԋ��@F���e�?�L���G���VFM��Ҭܝ�}��q^�Y����O�_]�@�FS�^�1��=�h� e|���XA�5ʜ���}�W��b�򟥙.�y{��D��1?�@�H��%pի^A'>:ʹ���#��c'���#��Y�m����D�~б�wJ�&d}�Ϩ#N�㻧��9Ώ��EΣ���[��\��BW��Bz'P�wp��|�����A��9�� ez^7�Μ!ec�"����"jw���eԐ�4�}% ^�$���Iv���k�N�Є�φ>TḎ�Y�<��-�M,�3���*<��a￞�N�4=�Dd"�+�Wu����N����RK�jiwIQ\�
):Ё�Б�CA��`��[�r8;~�̴7U]�]�<
Hd"3����~�7��F���PY��g~�5�����^'(�%���|\f>r�;��F��ٵ�؃������ƍ啙0(�3��E�tT��|p��܄�j�Z�����欢@k�>��K�dAF7�97�Y�%:�9�s^\ղU��4�~UvIzs#�J�\�Ŝ%ȩ���N.C8��Q^��n�H�!�y�T��T����>�\�ש`2<�O��p�NaF5<gP˜���Bx��YB҆5bfW(Ց|�2������JqԘ�G9(�+X���q�on��v���@8j��h��Y���D9����K�n�5<��� ��=���KQw�~�g�P���>���_�J�w�ys�C���������¾q�9��thң�BZJ�а���Es�3O?=��Ю9�������v���!7X�4��g�@f�q�
Up��۔�T�$�f+~��ÛG��E�ԟ�|rx���az����е�����ps�
uʴ����`�݂��|/�_�[�=�n�9L־�R�y���e{A��4�
��p��eD���@�kX	�\O��6 �u��x�eK��g�}p���I�ީ�S� ]��ͺd�.�v�L$*�|�6 �S����q��~�i/R&�U*\���(�]�ڰ�Q�EzWQ�a��XU斲9x����<f�~�;ޓ��k�4W�;
}��Q�@ćcM�0���q�.0E�d����x�{ɉ��X�W��M'�lT&|����bIS�F�@���B�{��n	�{;����~�j��:��QP(g�ؖ1^�����?I�q���B�������(�Mj�I!<��/R޹�F<�{7��34��FV=zγm{�`_�_��T(�y4�'�)-��Vc`�<��(h��||�<J�v���}ָd�+���V�|��y6M��12���K��t���D�6�Ñ�.�w�&٫B�������2���k�~��7O?s���Ք2vS8��N�Z�g1օQe������ʱ�g<XZ�|�H��o�Za�딭U��.�,,bU��ϋ�b=T��˾-�r�xZ�S�/�e�����9�LP�!�� 5�=z����r7W'���&Q2Z��w%��c0���~@���+�|�w�����؊Q�m�ok��a��5�0LyC�E*C�~ӭ���J
��r�)��2�$�����<<|�k_~����#�h����9:��e3���|>��zj�m�{��E t�w#�9h�u���9B�6���z�ס����h
� n�+�B�۷|���JD�1iZ��q��>�8YB}��z�ں�p>aK�ȏ�ﴷ�k��'>1<��8�d�N��7�
�[30�i��)�bv��	��	����g�6�D�0��+��`6n.�lf��Ƞ��ʶX�6�0/N3�z��N�
a�
�u���m;��h����3Dv lK�4�&�g��^��^�!s�*�� �������_|�TD�!M�#��/рR
~AǫT�z���&߭g�:����Ɉ��`�1�e��	�O�M�zJ����P���g����Шb�뢸�:�]���
�������ծ~�rk9�d4|�J�l��#�n�|�֍�)��"R1E�,PsI:c
j��B���(���T�Q��q4
<�3�w��wϺ�Iń��J�A�_�n_�o�li���x�ﱦMH�� �J��t�̲>w 8���dD�`#4�%���d�_���lG��dUqD���!9�d3�%������-�P]�+�5:u�2?xe��q��b�,�Y2��9��7��;�J�Q�������Y-���������}`�+G�x�܅���&��'T���� a\�Tt�����Xҵ���"X�
Z^�m�,2?k��Ŕ���Rj3&;��n�FS�k���y���B��@s�jcT��[�j�Tv�Λ����b��&
�v�n�y��Y�:	 �p�
^�2���o#x��K(n�d�~ X�鵌�H�1^�D n2.�
��m��qL�&���sl���Lk	b��SbrЗಥ��zVU��w�p4�=�y;^(FBp�põ�'��z�R�f�eeW;��D��gO=5�c`��]�]n��C�J�x��3\���ԗ�:��y�?�2��dZ�1�kF�w�ߨ���Tw��@@^<�@�&Bt�8k`e�@NOe�U�ч���[i~2	�ε9�J�1�)�E���]{����6�}f�XR#�E�hH����$(�mÆ�;�q��Ls�m�6��O�g���V�f��wNCT2_���:�����~�����v�\8��;�8��ȁJ��8)�-���Fֱ-P]ɩ��x��Ž`�9���v�LԮ����?�O������o��E��VX�R��u�^��8	㐙��~m�b;�8ѵ��N�6�^:���?{J%N��8ƇD.*�ԥ�`7�Uk5k�cAl4�����x�+�c*�x̍�)�����"-_���Ո�������c��:
@C[�R�����n���K~�d��D�M�)־O���W�'�s�N ڻ��ä����{]�������?�'����I�i��<z8)�*M� i�^X"Rr�H�%���FC "Ax��·���D���^�k��#���5�S�څdX��*.M׌ �̴�ёwV�po1#J����t��-Ґ����Ż�ш	~��`b8�	��c���ZF`E��}!W����*��y����������O~a��]E��vZn�ƑTy�8��c��c�LO5�.�Zd.L�F��|�,?�>�A��֭G� !ͬ���:������hZ�wPp�Ϋ�����-���9����L\{u���]�y�V�u��%S�� ,���<�==�
����رɌf,���&;u���2=���\��m�нvcs�����;0��6�Q�·��XכһË�[|ۮ�����B�0<�����*8S��<t�=A�����-��tj�7���Q���
����'�R�n�E��_�o��,!4�i��e���8��[�p�O����}��%4�O�g��M	�"��֕rk;e7dp�@�X��V�y3���xف�2C�;�N2�;b',#2���-��
��1^�.����E>I���G�f�3�{`���<�p���R�=i�����&�._�1�2�f�E�!���m�F�8sb�v�h�}�3,<�
����'-� E�$��%���S���H�yZ�J�>]R�w��,�w�<���c�7�G�W4����0~�$�~h�%9"�mi��3�#��g�J]{�f;�	�k4k���C�|���'2�I��ly���\�Q��m �M�1^8�:���@Hyq��To�%����v���2fU�c��_y���F:F��@8#d��w�U�8�DFDƔW�:�ڊQ�)�Liio�4FUƞុ��ٞ��ַ�4L!{dA���:c�\d�8�z�Dl:�N���=ua8��%�^��i�p|�u�wX �֜ ����\���I�C��5���`��a ���}�y�x�&޵W^QNX�Wk�c U�� c<��%}���T�<6��7��'�Rb:%�FX��`E��52'n!�
�x�>�V)t��#��c��g����8O�r���V ���ڮ�B�buǕm�p�Y��a�W�]B�[����r�2 �M��B��@�ZJ��.Ű_NW�8�(�p\]@Y��XRѸ`Y�Z�IQ�5t�Z���I2�y*aTr��1&$�H��ROE��PEzji7��c�	�����LT���*���ɥһ�n(U�{H�β�bh�\$�w�Y%���$��ң��;�����{ �J̑�'<��@덳�6Jx���/>��':���p@��L��c����<�[(�1=w�<�gsk޹á��Z�Ks'�o�O����P&W@�K���$gj�F&؂dM~x�K̽mu9*��fm��Lx�e�nBO�9A(�����Q�;i��O=1>�;�N� @��78\<wq���A��a��.�'�~{���� �x��&���?�������+.��P�� �׮��wT�����`�\�K�w�����.�bVb��]��9/�C?�r�!��Է���~+F^M���Qk��Ͻ/�}�	���n�\�^\&2a��1@��ɯ�5C���X\��W���x��'�O��F�ʯ���5$���2^�aۊU><K��Ǣ�w�1�r���Ly�}�:\Kw4D��h�pLꕪ����k����zԦL)�r����6l����%r�D%���s*<���#�t�����E�d �XP����%�>�����I;����s�u�ԃQ�-��q�F�0��1�R{"M�"x��0?T^,
�����لe��.�k��Zv0앫�e�c�{��ks\L���p~�f�G#?i�ȍ��yQ'٤T�~�B_��JGȵ�D��}���0�/��6�lɫWn([H"��nc�Nccl��[���y�%��Ƕ�3�_y�����~����]����O��-�լv7K靮CK1�:����G�g����%�W=��j)3܈�2g&zSkv	��X�z,*-��<
��+E^f��׫+�5��@	~����0���*-<צ*����}q+��-�w��+7lj�Oᚐ}ج�5��1zPe!+Nʤ�-�9�#,�}�;�U�� ~�0��M�bO�ڋ�* �27����{z߆�7n!�ņ��L�$��'��%�%�(9p{��@hNH�Bn�p��'�[��o�]�����fix����f�5��-��׹��P�T�8&H��&��~d�ZH�� 6��F��ܨ��Ry�kϽV��)���]#=�RƜ�E��8�Ǹ�0�D>�^�&=�ُ=2���X~�:��ɻc\|�+_��<�Z��?}8�i7ф�u��cPt�#��ɑ�|v� Q��\��ћ�����o}�ۑ�W�x�1I.�0j����S���!�'�}��j�I�$6�W_�FO�I�I�dSP�
��D���]��)(t��rҘ ]$� \ �\�r/ZFI���������[O�"s��x�����R0#�(]��6�%�*%���$��0��mp��a~(�Z&���m����L�Գ��c�i����Ch�{�0|�j#�]��Vx��m�)3E�`l��a:�:ߔ�73.�p҅��Iz�d�Mk�Y�}���+_��p�=D.\+J���FGa�)��x��)X����f���f���!�7�r�̕Ke5�{v���Ҵ*�W�qIu�i����!J�(��x�A�`q\�?y���+SLڢq)J�7�`��S�~t��_x�5�;�OS�_��
�{�H�q���A�J��ߢ����<t����_�����N����GLI�D�R+���Va�BC\��Bw�ּ���]	�߁)����V�H�\e(�u�P�z�-�%��6j������k��P��0P��!u^D�h;v����<�ތ��^��b�x�mg��o[ϓ�U�Z �p�\|�i��<�PP�}��A��,��Wv���q%zj�7xm�0,�}�ӟz���ގ���n������ �!�v��e=��-йN"ף�n��Zw�2���(�D��?��'��Ƶ!�BӒ�I��D�O�?I{�9�������c�/�s���f0�(�J�͒� z��5��;w���g?q�����c��L�hT>y5A�y�5��$�C2�|ψ�mČ�	'5A�o����3��N)�Jғ�������a�N�M��p���-�����(i��۷��ӱ'��m�6��l':aG6��pϮ�i.C���Umt���Ȯ~خ����p��ùc�������e�W�����D�KD����Fm���Yd�^��4��Nb�XC���x�x�[�a��m]�L��rr�s��w�v�&��m�u�p��2!b�ph�+�q�d1)Wm�l�a�2���B���N�m;�O<���ڊvZ~<iA���1��
\ov(u�w�X8��	��V��Pm���T*��> ���<W1,�s����hqJ[_ז�O��jW��Z�B�Z�[\���[ ���։bg��pΞL�9��5YND���^dYK�i�濍8����0��geLg�3u�J�ƾ��-��,/�(�
�Rk�jP�b�l����ޠ�dR9�翎����t��0֯��p�����c��.̽{շ��p��f�Qj�f	C۰���[�зl����w��k�w_~���$N��l�U���%˺<�0"��V�	aC����V�YU�1d�<�N�Ŵ�XQ����0��&w�P�D���Y]��,�p$ǳU	��뮞Q0h���X�c�k6���_ee�0W۾�H�(�2�.h�RD�x����u��M���~R���yE��uF6t�a�Q�	!O�2F�(EXM�W�����a�4t�/���V���=����?�j�
�OB|xI�7oC�/S:�)eb�jl�4k�1\�%����G<Be�2�q�W)�Zo�6vٻ�0���gO��0��8�P���?s��u8��:ӿ��"��9b�IGx����:����?L��4���u���9T��f4E��;,O�&�J�>5S�ݔ�P�.�͠�"%��o�'h�Ǟ>����/�J���TG�ݯ}�K���\��7a����Dr�S��.y�s���:�w�(���v;~�V�G��<����꼝�!r�OS����[#:�^�u؄C�_<�q\��=l���wE��!h�2[	��zܖ�i��� ��>i��:D Ԭ�� �ÆV����@�u�dp�`z�l����p׽���?:�ѷ^"C���f��nlD��(=uC�2ѻ7�S�,��,���TK|�}�a��WJ�0����N�MˈD�&UL��P��x��{���"�g�QD/fm��~���S���Q�c�#ytx�����������I����B ʠ�d�>f��+�%.��E�q��2�?�Iq�E�V$�A�L�)��.�D�b�G�3S����?]�k�EG��<��M$A�կ�9&�x�r�����YG���K��4Q�H��%�������=G)��ĝ�O���w�и����EW��w4K�3�R�{���x�{�|���G��� �InZe��ٽ��5Ž�s��y�wֲǨ�U_�U*��
�o�R�ň�*KH
ei
GJ�D���X�k�O���/�����ԮL��S�{��5u��nk3�͚�4��U����_6��\�2o��x��c������q]R�������{e���+�&-��9��q�ׄ��"*k����F�v�4��$�|彄�S�Ns׎�����?��%C~v�j�������h8r�����(�q)<���F��/������<�|�&$SX��U����CI���7��h�-v��>�9��%r�o�x������?{f��W??�s�]����3m�̋��?���{�Mr���m*«E5���F��<i����>�&m�a+�b��ukC�RBB�g��~��/��}����cg��|c����[�;�ޢ�����W py �>�����W_(o^��n1 rw_@�|���"U ۩8x���<j�(&s�7{!mI���xſ%;O�9�!(-+��)n�u��%5q���VR0�8�aX���gO �˽tB۽�s�Ϟ��"E#�����4�y��=l=��%h)��"0�I|��6�a��l�pN/�J �.�3Ģ"&à� s������Sy�t�.�|�*��0ȯ��H׼�(%"oi�J�A���?�2�3@�%�{����Ç 7�X��p���˴Q��P�����B���V��R��
{(���J�X�1����#�-M�W":������҅k2�7j�g��&��Y����;y�"��e�2���Bq���q����uu�5YX��B�wR1�W�YƉ�B���֩4��$ұ�$sc�@இ��ި�u�r�Qƹ��po��3�k�Þ��U�{wm9���?�������;R$�ۍ�̏W~���jG+,�{_�e�zy�	�6����j�r�}Y�1ݬ7Uv�����	(��[H���:)p
<g�iҚ$���Gf57C�k^S�#��0x���!G���1�sݖ	
��M<��w�G�K�Q/z�3�M?��K ��s�3�`a#�3�����R:��!#��g~��_���XƽlD��s��!�;���c�B*��`F�z�ό�}�ci}zLj[!ZٶmԔ/�` P��a~^y����{� ~�S�/r���QH�ڥ�=w�B����e���,�kMX>2\:׳^'c��/~ƶϣ$ls�n8����Os�i�f�9_��?�좘��⪬�{���m�7"���'�D���V6�]��)
~�o�wf8z���*���^#n�&#�҅m^�������/e�����9X�^�zI7���������;qb8��4as�l>v��������K��z��$��e	͆mZ2N��3��,��
}��<9U{ �~�V)�5d��z����CQ=���o��o�?�di�{�^�#"��h��q=Jr��q���p��� �����KKj�~?��ہ�4�,�0��I���oL.�ߊـ���(3��NT(3S+�V�W�֬�:�k�&]���#n�WSf��{�H@�и=����/y��̺`�v����/�w�F(�]#L����w��%�5�c0r��,�*�5J�%E�]k�Y����-T$$����)�O���;�W��5Gc�	o6�jL?)O=?qz����_o
=NA��0���{�y��1Z��]���%�)P��a��ņ���c5O^CZ,�<^��������ڰ�ͮ��1�x�#%:A��߁�2�w�㱇�g�x��g����I9U<���s���p���5�Y�a�Ҋo���D(�n�D��k��c-���dE�w-A��J�N��1�7c���OJ�������]&e9�)˙��[���4�n��zфI�,m���4�1) �qC�l�����[u��C�}<�$Q���<%B��]���ᓟ�ܰ�/�ia�(�ؓ��m��wJ!k谾Ma� x'a�250C�Q�b:��Q���h`9��۷w �߆�� ��V����7�%�l�T���xQ��̅^ ?|  �^ji׏�Y3[���nS+~c;��_L����K�W�f��"͘=���A���Ͻ@TPʒ�%Qė.�^z���9�O~�b�,��$�n����a����Ry�z+ˤ�Zܤl7?Í^�(4��Q��3y�UD��_��%���w �}XU��n�p���p�<쮝	�26���/e
]�"FM����?:a�}��í7iȂR���Y���O���V����.,�N����6��OS븧P؋\�d9r�/��fHl�&��1���o��'��U���W/�?>9��֫ÛP��Zw=`3p$   IDAT ��sg�W@L\���שHI����GR�=�(q�e�`]�f�ӻvS�G�|����%j�W��H� <�&�c3F�QV+{�4\lz�r2�y�.\EIHH���Ű�J/_��h_h��C���-Q�D����s�6
�:|h_�yS����ktE\�f��zɇ�������p�,� ��n�<���N?���kF}�$ʽC�h�"v���E\E����Q(<wu�U���uu�a1�WO��,��~N� �}����!�}#�E��T��	qT���~���!�Ns�]$�˂��֭���~!��됏S�O>{���1���Dy��`Xo�`o��L����رuәO=y���_�z��.�!��M�#��4��^�9*:J��p��5�\u-�����%���Եqr����"����a�u��z+�o;1L��p�g4��k�߷�f���-]��2��ɵ&/�񻐚�C�O�y����� ;��#��	"�)�w�>IXj�*���>�R(���X��'�dNQ����o��ɒ���N���ƾup�I2�	J�P@v���[zQ��L���.f��P$S!�XG�}3 .�Ֆ��x��@D:G3����{(���Ո9�iǦL��s�]��~�>,���_��㝆8��u�'��ƅ�����2���w89P�E�^<:�-� d����C�_���c� d���7�S���E�4x[�z^JŁB5kb�e��hS	�9Q����zs�+�G���-�3�#�-s��= �1<�1�jv�}�5��1@;��N�B�(�����e8z�I��g>�����4�X�i��.�X��g�NtK��.�t�ˆ��v������7|�k_L�ȵ�X�D��(����}ï}�K)ۊp��ˍ�,aI�3�x�u�FB4��W>W���L�<p�R�Y�SD{6�ʄ�%@?��7���^��v�wΞ$�����o�9n�zy�:�r����/
C9Yb%��{F�]��F��Vߔ���м��i���>o��=f��b�S��r^:OKң�R�~6��K��$G|S�ԩ3�(cؐ�غ�ѫk���]�DK� ����LYY����)y�#������@Ύ͕5�S��5P
�=�w pS�~4>�m��y0ߡ��s�Oc�})!��}s�^�ޔ��9�������e"(�]t�څ�2GqF��LR\`�X!�*J<ӚXc�	�vK՛C�!Me�v
�[�/Wqn�
vv�3�s���M�J���u^�;����gXf+�֑��=w���o��KO3�����.�{X�gnҸ+�rU�ٔp�[��n�}}1�3�e��Ϧ�!%[��RSC�y�Y 5�D��S7)*�M�a�B�V`�5���$A1��U��Psj^��z��	��Pg�!a�(�Q	]�Ra�s�E&)��kž�\��a��|�S�L��	���g6�?��%����5�^sjfʜ��b�n�粘Y�q��w3j
~�I��aa-o�x%l�=�^�u�� �}O����E��^�
��;�E �Ea	tQ�o�]��Ӥe���xtR��g���ߖ��Ǐ#�~Iu�e�C=0a���}P�.�+�3������a���a�P�8�&���.��>�3 �g�tv�4���p�R���j���kU�W���/��ʩ7�o��!]C��q� �	� ���D�e4�"BO�G�<$�˩`@^~�C� ˗��Z��zJw2����w(���A"�|�u�*,p׮<�;%Y�� �nP5p�p��y� z�(3���݈�߶g˰��^<�}H�5=4�{��ݤCLsT�9덥��B�S��gݱ\E� �S��;�4v 㬰V}t�f�T�Ft,s����MM��=�=�%�ћuo�r(ίwm�Pǆz�1�܂��_!��@����$�	W�%�(�%���3�g�\�S^�v{=�G6o @�r���m���ڿ��3���0����t���*��|��!�q�L�[6���h��S^KU�p|tye�j�-9��+�ޝ�ȟ�%-�V��U)8���X��w�=����������Ż�h)��$�M���X�R `S���L�'0�&Ѩ�qN���X��A�}׃�Ҏ��bL�MCvc��N���S�S4�_!�b.�ֳ�_�^�^>j*���=OdpE��sy����y�����f��q�,��&����@�+���"$��e���������K�}a~��tr��D���圜�!P�pܧ�\�Mq����QZ�Vv&����Z}��t3զ���B^�ҵ���Q����5�n�W���lFØf[��	[ī͢�+��r(�(v�=>7)�Ǧ4��
�i��(�4��#xƳt)CH�=�k7�bl�M�N����>�ȣåk��}`-�C�[ o�^PP�Bɰ_Rd�^��Ԯ�s[��קj��
l�jyF�-(_o���Fw/{������\��z��Ȍ>�ƶ���ˌ'������ߊ�sp��t���������!�R��?}щ��aɟ�y����>?������3������C����jQ�C�UJ�n�'��8ky����k��x��w��� tS2�]��%�QV�����MWs��i��g����)B�A�kt��o΂!=�e~0RTl
s�3�߲�������w�G�/3^��F]�g!I�a��O�1���&Dy�����w�	���!L��庶�-MX�ߵ-k�P���}ix���׿��a���Q�B�v#,),�~	ı����qu�J����q�4M�,ˤ'+�y#&��W�g�̏�����5��^M��p�ܠ���w��4�n(︩:�M>{։Խ�B�y+9ߔ�aL�/ʧN�IҟbR�s���xQR"��h�}Ɬ�N�$��=��m{��)<ދ쩭܇��}�ꆅ��so�Э��쥌����Pi�5y�z��H9A�+�%@EdD�Q��v��.��&K.���,H�y.I���*4ܛ���'�޿���ZJ%����!�Iw9&�.&� �OR�'���H�T�:�K�j�rxb �4�Jvi�o�Ny��?���1_�B0I��"'�UvIQ=�a9�v.^G��&G⸭��������:y�FiН���:�� ��,�u B7Q���kM0�����dB����+� D����/�f����Ͼ����჻�ڶe���k����|�Y�Y�|1¬��K-��b������ب%Y?���:(��� Q5 �lY��Zzx��&W�V#_%�&+5��ZB������ZZ�*�7L�MKī�׸������*-QAx	>��3C��~�)�0��g�ҙ��~�7~}��'?3�M���?�%߷��������JjcJE�D�δIHVȣj�+�h4�'�rB�MIHf7��G�=\V�r�9�/�vlx�$%*ze�ъ� �=�����*m�w?m Q�����
'u��[�m5w��-��?��?E!��瓠��s�F�ʹ�\�Ar��J��V�[�.G���K��g#@�c����pe�S-�IP�y��Q8(W9�7m߭X�ב��G*@C�x 8m�⨨8�"��fg�ۆ-c`�*�OJy����U��u�~���a֓En���s|v�I#E�k��/�>�w���O=	z{wJ�ާ�t�70�j�v&����t[�V��}d��Pqz��yǍk�*aRk�mt��·���h��}O�a���s�'IL/�4�SY�G�ʬ��84U��X���]�z�f����w^SI�$�o%��G]宁gT�p�5"H�C��Q,s�c���)����¥�wm�wH�=GD�hɲ�!]a�K�G��rͨ�
x�fOڹ�u;Ѕ�^/?.Cɢ.��L<�R�Պ�=�_JFm���w~�H�|���F���N�:����L}P�R*H��%]!�`�E{V�FS�Yl	����j�UT��=�h���Q=�F��%���á8��Ð�<0m���^���%o���I���*�C�)��͒�g����ȣ����~]����ggΜ9���G��w�;��0���[A�'���2�^��K��O�����B��ҁ����7���uǮ}����z��g��^��JE^�Qy�U��|�ۮ��s��*�Z�Q��FmSb�TyQF�Ik��
�z/a�&L�'Ne�{��Q���d�T����"�L�eI��9���T�CKڒk�> ������"��V��!*�x��	��+�_����-�YM^}����?J���h��y/��-��Q�������ס ��]��6�1�d����9���}�<)0�9~��9(IסP���?��0�n�<���	�ʾ�Si�zk�Z&��EU0�P�i�r���pZ?��(z�P����������ީ��׶�'��硿�x��mx��8��MԺZe�o��@޴��-���XBG���ـr���
��J9�ETt��4����+p�V����e6��D��M-���eD),���M������TET�W�[Ě(�ϜuX�4�l\=��:���(QQ�z��p,�����~j��ٿ��9؆kW�%�:0L�x�_�b��q����DE-�E%������L.�֏�[�KC���3q�~bx
�)��\g�T
�5���������fW!������*�5n��?��Ea���q�:��Q�����^��d���*j7�n��+�y��S�� ��`P��|;������4����5�*��!KX�w �`����FH��f
$*�~��5���ipV�ըb��x�h$��M@a�A������8�.]:�:�+���g�Rr
 �c��O�%2v  _��0)�2�zym�%�#s_t��=ȝ�G�4�w��?���vqn�I�H�5m~��M��cvX�YX98��!qg?�H�2��o����O������M�lCf���ʱHxK�P���&�5?~bx�w��w��K����������^=1�B��ށ�a-��)�Z*Z��a�����^eg��?��|���6���\ˢ:�94=|Q%�O+�𼻕��Y����
���h��i���q���"�=�0*h�ɍ��k�(�<��@�u���\�}0�݆bs���[g��t��3i5-p9�}��7�W`esL��'$��1��иz5�p	�4˝y��l�QR�6��1��=�Ǣ^�l�����s_���Ly���)�E��� ol�4�����x&֏?�t��{���zX�.&�.��yʵ.#D�?9��fx�╋x�(h��' SQ ���+�ߢ��p�#�u����y��e:�� hs
��4h�M�\_�Z�.�i�L	Hm���lԧv7+p���x����5I� ���1s�G��*�W"6��XVS�<�&�r��v��t�T�(`1����=8C��0s�u�BL��Hs##��ٍ�l� pr�|pRx����N����u`�v��`=;OZ�����gZZ:&�M[��;aw5Uc%^��DՃ˘�xd�a=�Z7�Ʃ�� #�i��{ډ�d4�j	����S�yH�����ϕ���A������:ɕl�Xe�7b�x�brR�ǜz�@����#�]Z����C��F,����AX�~����X�{Ħ*0ĭ���M{$F�n*:�C�y⢦�ϖ�o���eZ]q�#�zİ��+G��%V��҈Q�z��ƹi}x�H�87����V`��#�脚��]�V�()������O�E>�qSUE���p�)���[�Uhf�t#6���w�t�4�j.a8�h���q�5M#{�Ƹ��F��y���qw��H��$N���˟�Kߓ0e�Ͳa����`���8�m�9�1��իsc����?��//8rd�ʆ7�����%�'j�Fb*�lH^�Xÿ.�"7���
�<(���КMu��X����aǛ��G�'��煐�Nu%>�@4o$�X�IՁ
݋�]��}�@d�ғ)O.����rb��K��i*����9?=<3Ӈ�SL㍢;�%:�i���کKo�{�@���}��a=1���ئ����3W��|����
$#�=fd�KƘc/�/�kq�5�����|��+�P2����I��N��)�Z0��G����pmx���ၻ��m�$jq�w��'��m�zʓ�06�K?���������[�3��w8��α�c��BJ�^}���_���߰$��U?`Z�{�K��?2����õö}���H�_���w2,���7�d׳�Ab�	�rME��g���6{|�0��+��(�|�<k��݆��`�`|�"ѕ�aˆ�Y�z{��	�TҘ|;��;{)���h������g �%-�yB�7�X&0���ݧ��vq}�v�Q������瀢���(^���r7�n��u眧v<�Fj]��.�x��&��S
?u�*Q[`�	(�s)��1����Cc"���@�4)����^�͂�gM�g�R#ʗ��� F������MR����i�k�Gc4��8�6j�ǝK�
�v�(6s�+�Z1�&0� ^Z9Ri�n�t9e>ηQ�	��@	n���y5ũ�X�f����u oL�D���c�TT������\C���M�D�8��K�Vj)<(�q��,F��=����OzcF��w��8K:�{��S�v�؅��X���?�1�	쿆���7�:B�[!��6Ǚ��@�h#r`'�4n�y�ell�BX1��:�ە��#�ޑ
�|��+W�����Fk�u%�7S�g�k�;�e�*���� 	�]�����7�?�%8T�0E��WCI[~��S!ބA̾Ֆ��a��vQ�6��@������+x|7�ӕxb'<ͩc��*j�i��v��c\�7*� ��ZK���r��-����٧ W9S�f�i�T�����)���QɋEl���v���k4do����/,�0�����-���K����^��PSl����K�\AP��K%J����>4R�6Jƭ]C$v��\���K�;��<�0��9�W��?ǂS`���\`.��֓��G#���
�/_��'oE�l ʰ9\C���6�w������@���Ȟ8y�\�g��g��ǟ��ߠ��������<ш�B�d�̟�Ռ.g_��g�3s?�N`<Qs���%m+V�-�6?v7��6R�Gͮw&�����dK�k0�8�m�����9kՈ��@ ��7�P�J����W>�E�4��R�r�{�H>r���[�AD� �8��:x/=�w�N���c�""s�����^j���KxY���R�!	ھ��1<zs�̉{,���3o;�4��GaSa��p�����)e����*|u�"@*{�k<��V� �|WJ�*/<@�9a�I2њ2�Y*oհX-Em�<8� �v�u��=])�� ����o&q{����}�Mj�E)���-\���D�d�xp��H�m��|(��ua�o$"b�}�X��˓��T��.����īL��z��v����k�y-2
�@���w�h]_ZEg�W�?^�W,��{vo�[��ƞ/�k97��7���p1{v#�� �i������x��?ל�er=�Y���\�r��D0����{v�[7|���sL���~���W�&�^� $�ug?�H�~�ԩ#'O�|�H	Z�g�}�k�\�n�s�K�IJȓk�6�6��<����+ִ���ʭ�{�&- Il�EBD�(�śsxy�@\'$R�&
��XS=��[���%c�;�E��$��4p�������Z�s4���5OKp�x)��WAf��\��2��xM��n�̳�F�e�bU'�[�\n��Jql7�����J��S���KM`� �������b�����
Ԧs4�0�+�ױ�4̰�5�цʧ��yB���T��Rꞡs��Z�]���F�	9�Ζ\��*�m;���_^y��S?�MZ6 �[��(3�&ϼg��?98xdx��W��������tl��?�6ㇵ/�6^��
䓟�7T�������_O?�<as��o��0�#�>1<�'i��8y��a;(�6Rw����a�#wSK|	0�ld֒@E�!;q*�Xza���[���0{~�Da3uT���0��4Ѡ�z�T��A��r�m���f=���qHtf@J��:���������$o�>�Y�BD��W_�P;9���Cۜ(��}[��3��/���0|�;�a��°�mx��	��a�!ް�3_��D�l����w�f ���xSU
֍��\E)��P�p�bK��Rajy��i���h�0��|V��2"��*R{�4���u=K�E9�Vl$Ǡ p����{7ǟ4� ���@���gs0�V���-�#�jS�4�߫&+�����C������f�=�j�ltG^�TwW���N��:�:޺���&��#�+�z)�b�@)p�aq"�`�h�YQ^�L�t�\U��C��~§|��$��6�zj�@�D��b���F)�ܽ�����lX�:<��Z�!Z�x-"gM�1:u�-ڙ�;{8<�1rɮxa��K��O}���U��t�A:�8��ݘ�ٹ#��������I+��O�}�cOgE�)�Z��0���J��^�Y�r,���az�aRy��� +ih��VN/�I�h^,����"�3�ۻy�N�3
������R.D�,�V��Z�a��0y����}I�����uLM��ܼ%��dֹ�mEY��1��8�}��{�2���d*��e�I,/���?<>~/����1/�cv��"u'���x}w�;�H��l����*�1��o��2<��e�ȥ����+Ϧn �[�y��+��� ����1x�7 �D����Bk	��m�l�R��r�E޿�k�@�ior}[�������={@�~Э�
vD ڿy���ã�?>9�o�s��e�;�?�$u�0�!�o���۱��Or�7�_v���������!D:#rnu��AY��-AZ�^f��1�)VÖM�v1�i̼9�����q�(�~�K�n����7o�����H��F��9�3' *�t��E�V�` �9Ble{��n7���/��E~�����X�4<���ý�>8��|��&
�j{��U�SC��S^���U�rd?VɢUU3o�Jo�P}�k�ʍf��C,½W������(I!�et�Q)�2���kz�r�e-
�2����x�B�=L���R�֪�M}z����[Qyxe�Z���g��c���g�Lm�5�%H5��>+N�D%�3�-�]�'�v���-���G1W�M��y���0������.J�v#��,�������h֚����U�2�6�W���z�y�Y���*'� �`�H��{�6�� �(s�M3���t�#�~��0	6F#6��ѱ�TZ�N�Bރ���r��q���C��Ko��2|�3������9�L:�$2�f����8�n�o}�[��A�_^��X��(�<�z��E��z�*$�Hy�.P���Sh{�fO�AY� ]���p�����V��`^���������˽B=	�!X�B�)�E�P�T1�L&����k�
d��L�*2�AJ���O��|����P����+�����������p����ٓ�-x]��W����_{��h��H�^��vj���z�8��`	oE=��iȴo �6�N����}�;�^���8V˝�97��R�FTz��8�����\)1���P���z��P�2���%	ḗ6��Y�v�x���C��#��M���`���u�@z��!��/�K�,?F�$?�n��'?����o|*�Y��]��3��=���{`�]8�#Q���?(_���(��n&���YG�b���%X<#��#mL�5E��%������4�'�ӷY��>V���w_}���9|��?�`r�(�R Nӡk����
-�|����oE%h��,|��vh{�8�~#8B�{ȋ�ݵ���ѩ�T=l�0(^�����u1AM�}�e� ��جE���T�,'R����*hhS� Ī�-u{��+��27�?Rѝ~��ձ�J�E	������f3:����X~�?z�^#@iS�x�[���|��gYثƇ׬7��ZU���O'R5�an%�a�u	 �����5��,Է��������:�L��H����R�f$�Vz�f�^]s9�e|�,f�IZ���?P�>͞�c{B=�����i}G��|ט��|-)PC�R�{������O�����wŎi�@-6�5��/��c�� HSeas�%��H����s���N0<S�dY'���8F�E��]���q
���an��.��Օ�����X-ބ�0�W�2�c���7gABzq�&�{�����^�E�j��ўoʂ^^�:���K-��!��Mc���Z�|$H�\��t&,����Vw��b�1S�{���)B��Kt�EX1NE6��K՘(�H:�����A��n�@�w��+�Gu#I����w���g>���y��~���D���&����B�*u=����e�T�8C>d��K�'��	,L��j�R���o�)$���a77�|�O����#�d3�]�}�ʟ�ٟ������2��K���>����j�5潯���M���µkW�9���!�Y��h��2
A:;Pdy� ����Sǆ�}�Gx��0���W.۶n8����ǿ ��hޛ��q�TX.�H��C���D�G��Q�+��9��� ��f�Vk�Qҹ��%�#�b+�I;�ɰ%"�҅�Ʌˌ���ު�����t�z��qx��'� �w�J_n���ٽ{���{�)L��fTqæ��&hUJ��Ш�DK�Y:��Z+�כ��@���_<|�Q:f��JPy"����p�K6�_)��0�5���������%؉<p6o��%����׹���!�p�3KM0�
��k7:���5�P�i�,c��uվ�7)*����J*+8��Kz����M��S���oʥ���rhL�.�
/z�ɨ����tS����Ys��ʊJ��/��U������X���rn�^���Y9���m���6�/�sߛL��4 ����-��m�L�D�؍1���dL�/sź��E�i��%��sϾ0\C�ݼ��)t�f��p��W�N��N�_�6�z�v�ǲ�m�RT%8F��d1
@Z���N@�C��<��
*��+ ��Ʋ+�,s8�Fe��u��֠��{���oi-������ ���cK�e�s0;�U%r��Y~�c���wNʞ�/��]��>�$�,Z)jK7�����!��%d���B���=Zk!2� {��
�K}^��#�w��1�ع��!�	��M0�i[}�����M�]�=�֞3ɷek��\��yqL�k�֏{�1s6�X/��(=)����T�?�;~��� �.�^sk<�����k����o���5����4���8\<w6�Y9����lۼ5���#o����֛o�}�I�~^�Y��s���j���O��?pee��7��~w���ߢ3���e�jo�;O����ې�,P�n¾I�t㪍����B�>s�Fi$9��(@ْ���Y(ry��D) Tѐ��*V	N�>}��ik���9@�=utx���Y3c���q�rܟ��'ׇg�{
��/�u���}e�C��}򙆹w���ߑ������F@u�]GH�Ѓe����
Wp�X�~��D>V�,���V�.�=�V)o#h��ve�Asz�v��;.#���VO^!�R��5�*�ev���s�*�|��#Q���s.��7!	�\B�ݨ(@^u?sYW)��H��}����*��[C�;^�?`(;2�Ej�ZY�)����Zk`3�cٚ _SEa�[uh<�^y��̀Lz�jR_	���l�x����ｵcf+^4�b�T��x��Jw6E�j�)"�!��I���H���%�[M!��A����tu�PQ�p�P��"�_:2���@�ۺ��-�jkc�'�}FD�M4��Ϩ��1��硳�& )8�l�rΆn4�2#�P9�� +����f���N|�A�����Z����5�/����c�G��[�3*�l(�"�<�c�Q��Z��
�y���'y,ȐW@y�����}gq�x�89�5̃Z c��+��j�+�'�h9�E7u���&��J�S��&�R�\�B�?s��qΛ�H�
;a�e�c�Q<����rs�Q�H�����Q&��L��N���K����*��&L��#,j.���n�S;�l޼���թ����+y��dx���1<d�CQH�b�����!1c�I%`�E�X����N��B�C䌽��Z�������{÷��� ��_�,�:����_f>��O������n�Ќ.M��frFx&�	9�,L���I}�JV(����*:�.c`w��>;�I[����E*�;
�G�`6`�,Q
D=8�w��i �����[a�ӈڈ�mH��Gxax�����H�M$������/h�r����ch�K���q��hﺧ�ʹ��;�M���C���<����:aޏ�ջ'T/7�)�
o��,�z��)k��O/��V�r÷���8���{��&/95�A����;��W�t�[�=|K#Ğp,�2�3�E�����lޏ�װ(��I2����$q,�0��≶��;��퐳�Vz6{�sf})�HU�Q��i�����;VT�)���zV�r_�m�5�|�xД{��\�9Y�;�-��5�qͦ����;�&]͘�Ik��X;wFO=��:	5��Ҡ��3���m���b�)\	���II�������|������#�.qx,��{`��B�����KȆ;����:�mP�=�ܬج�Z�k��B(�4���\f���i�g�i1Sn3��>�^�z@tn<��aF�{Nar���u�.��/ٸAʰW+'gs�F��1&��C�TaC�n�p6:��3.���L���~�B�s�Bh�ܪD1��$O�aC�J*f���Sm�״���	N�����`�������-'H�h�H�Q��ڴe;�Q6䖝��\;6�d�����9�$'���(�|����"d��$5�����e<���Y���s�s�����}������ӄ�(���tnnx��W	�����?��&�.ԯ��?~ix�w�	O������ �J�|�`��!�|��������ȼ�2������o/F�Eh���	<ѷQ���|���a?!�'{hx	p޷��x���x}�k_^��������!�g�PP_�i/TJD�lx��Ѵ��A��<(�D�<���f7�Z�y�҄U�;�����`>�z���+�0?����kg0�v ,���޿�����-�?Ex��a=�7o�J�����׿}lx��3����IJ��1���t#��2|��-��CJv� �{�!j��ʺ����l�z/�*0��.�i��h^���+҄�y�g]���\F��>�e*]�����U�w�v���qy��m��=�����_���0��ɽ��!��iŔX��*�g�L�I�|T�:��ngDo��*��,���cO(7LA ����L�-����
�7���2�43Ҡa�do5�X9���*>����.��1�#�w*�����c�Δ�
���(��(y�x�S�����u#/�H���;1u'�U@�6ne,6���}̋��$goy���D�\"�IO{֛�8�K:v1�����l	`�[C�����0;�%%��|N���VB���q
n#�"|�ee��T��s��n�o�4N��}�(,d�BA��B��7�?�gΖ�h���.��$Jgލi�**�S�;fH>��*QQI���JS����W�6�һ�s�� �;6Ӱ�~��� ��t�O�}�� ��S���5"B���{��d�����e1�6�/�{9�
T�?���҇��`Y����G���I8�}(˴���]�	y]�4����6}Y���~��5R��y�gZ�][�O�gi7��I�5��e����zp���'O�<�}��D�~�� ~aN����hs�h|��:��y����W>�	�{�ϟ~*|��P��C�z�_Ʃo~����3�������׿J��j��×�u�t���OS�n��[i�"���+��'ՠ�oC��v#\�n�����*S�V��a)�F%oEr;�i11ů��j���[i�J
��U�C����p��4�/,��8�>>ǜ\w�P<��~�3��=BNCQ��&�o��:q����/_^{��1;���'>9L������<|���&�����;��u\
�E#��ඡ
�B�F}k��؁m	Is/��C�*����[Ei刏B�WT*Qb�%f�h�4��Ϻ���<Vg��A��s>��5�G��{�}��lͻMN8�2؋;��ι~�f� 4��g�P�h��K>W��*(�t���7i�Sv��M��F���N�<Vs��f�M۽.�ȋ�߲���@v]���`��C���QR^�X������|�S䵷��x�Ց��YS���4�@�f�HsD�^y�d�-�����L�����h�w�>�޿�)xD�� Yv�ȡ#�,)7���J�-r0k���N��4沝��TJ�7��!c1ޗX��Ww�_�<�͔*�*K��E�%����OV�ц��#
�l#��� T�#��ɔ�n�H+(���n�e.�+������ G�T
� @1dS)�)������>���r��/ek���@����sj&o���j��-/�+��f(�Rи`��=�^�S�1�W��|��7J�f����8�T�#$~�6���D� ��qi�� �&����l�#�����(#�
^�)MKhl�1��!���o=;\#ל|j�w�xyç8fRֹ��'G�k�]X�[�>�uj6�ܰs���O>1|	������?��!���DAI�aLۗ�/������~��p󔶐���&�ٳ{/����>7�_��=�Cy	P�b�����q��˛f���n<���&�vָ���;����Nb�RY�~�#@��2r��a����G�R��'��/��
Į\h~FzW��G#'Dl4H+�A8rÖ|r�6S9����OcpyXtDS�x5���g]v���9�{�$nM�.��⇯s�*�'�)��uHe�Q�{��k��U1XX��x<ɋ�'#�(J�r��i.�[\��*$^{�{�U;^��]ڌ|:mu�m�T5D�S�֍Võ�=��yG�w��=���=g��yM#eP=T_)����~-Ui*K�vUBW�#?����9�ԭY0 �{����M���B/���D�zrƽ����7*��������7e��bP�0�qf���B�B�!�,-á��4���Lc�-��C�	\
�<4�����}��
��K�c���apY�D�^���w��Y�^m>36�9u�ʹ?~�RFJqSx��o"%6�!2������;����f��~�s7Zk[�j���4�,���8F�7:v'�/Ys��8]@JyS��<�Q�,H�ۿ�\����YңY���&r�	����#
���|�£�}��*��*@DJk!ZRȤd,Q�*�����"�'}�4MHT�+��ޒ�Mo�����: �;Գ��%0Ap����m�o���g|���BWc�R2r��?�5����ʖ�J��F�)ޣ���Ux<�8�G˻��}
�Ǉ�߆}o��"�ۻq���?5��'p��/��^y�h��\Ǥ��`� g-����5������_�M��p��O<����3/����3̓�Dy�dӪ8=���'?	(�������?��H4�x!`$n��/|���D��=��*_�	M��pFs����/�a����K0I���W^O��M;Q�S}���g��k�` vC�b�{�3�=��%��5� 4Ȱ}b|��]���r�c^���KYPи�`�\��B�"@� �m���z��.5c���??{��̰�0u�m��EVKM��FoX� ��
^�x�唧}�49������%l�;%�$��t"p�Kaj����Z�5�Df�hzs�����uݮ庽�^:V��jD�y��1���d�,�����X�ʯW��iT�=z�Q�1�/e_���纛U ]k�2���y}�d��yN��x�8˒�P޾{@�Jq4vY�8fW��j'�˪E��;x]���^?+���U��)�f@���Hd�7�(wٝ��3��������1��ˤ����CN�〔�km��,RW�� ���k 8�,�vd�:��r�W�4�#����W��)�$���� �F�ڏa�)p3�8V�6�x�-	p<��`F6���#ֲ�&��r�0rk¹���|�Q
�M��G?��,V�����V������hÅ���L�^,P�`��[���e�*`��L�Yeq��ꐕ\Yl=�[�7�Z>���d��]�]�v��+��9W����dfj��Ά�����+^�m���zhOm����%�o���{Q�����E�{}��a��yJƮ\�?4�`�l��U W�k*48�V:��M\������������_�2�.e���M	́X�n[�n׻+����<C�nF1S p;������O}�zqx���	�/��~����ç7a�+ઑ��6 d�]�0���!ex� �Js������n���3���dO����I��v��4���/����{��<���O�����!B�[	G?��G�9Q�O���[���7Ŕ/I��Z�f�J@ #Q[��Py�bD��۴�
bY0d��.g]��׻��-�}���[�����rO�5{�G��q�r�p��Aal��M�T�N�e2!�Jr$�IL�z�0�����9TZ�,��d�3��V�(�W!������cG��1c�q��{di�3����{޻ל�ptO�i���,t]9�Z �|נ͌T()��{�}?�Q�v���[}��GB���u��~n��̬ܽ^2�o�T;��%ru�a���e��5I���ܱ�h5*B�f�ٟ��ȇ82��Onwɓ�1e�t�\T�)�j���N(as{k�ȫ�p�}�O��g��_��p>�����0$V����0��j!{�X�l������ѵ4��l�Ȳ4���D���HS~��|��oڴ%�OβOg!O�M��F�w�$ߟ+.���H6���c���W�PɞCc�CcD�����������O6�8���LW�[��^��Rh%>|��|�Mn��6�����,�Iȭ�a�V*2�t��j�$����vd��^�Ql��h���]K'�ڣ�G�l����YU�����{n��[��p:d��*^Zh�����ߞ�����Kn�����S�~�l,�m�9�P6���L�?�ϦәD�o �d*ہ}��Ki�x/dQ(\��>K����DT�D��C�x'�5������}L�j?I����?�]� ��A�g�9��w�����Hd��2�Ԡ���2˲L�m��ݽ�����y>��!����!����r6�������N����	�x�)�H8�p�e괏2{���� h��Ƒ������0 'FJ�4R!�ܭ�w�a|(f�"^$�0K� [)�R���R%�#�L�b�p�"Q�׋���K/?p���y-��R�o+�����m�bZ~ @rT�����@�8;3I���x��`/��s�ɿ�]V�)�*]�4Ft����,&�b/C�{��Z+=��7Z�֑𣯅��s5�|������Y�^��D� �w�=�<�����n���8J��TB�_3Ҙ�nxS@�K�A� U[ Mf�H��	1)�,�P���c��M���W��F�E�P��H�e��oFs�[i�9�U�ՅLˑGV4i��r%���#�6�tM���/�f
f��4ڀ@i���_�Ѽ-�YZ��(�#d{��B`��d7�S��b��j�{��H�á|-�/FZ��rz��=�E�;���ߊ�p�Tur���HlAm).����;�q�y���>��F(�� d�<�nE�NK�Fk
=��'Xko���,e*r�Z�m��"����Je�w�����nm�x��{��L��4�&a��ΑQ�k+�_ @���,���r��3�	>�X��pC�Z�uWX~U���إ���W��A���,��a@��S�w~�\��q+=�������:!Ϋ�$b�Bmۻm�����@���8�>��SO��ng�(y�8\#�o�7g��T���WX��l�}Ζ��_&��kJ�1P�\�����F\��:(d�%�sM����kxBzG��������S����y3s��~���(�z�P3�5��o�Σ�o��������}�5�(p�+c�o bq�<HN��T��z	��e+FK�֣c3߆��θ����'�u�R�f*E�*ذs��fH"T��д�sK���V��9Zs�\]�^IB�K���~���Хh4����6���y-�N��A�G��h�7BT@�y��M�����4���AџV�Tŉж�ӛ�Q�Q��k�k͌���1��Z��w�(���W��AM��y���8V3 z���1G[�f�DqW� �y���M��g��k-������F/4g!�Z�q>}R���k��M��Wࠨ5]�-ͷ��w�D��0���.ӡL�Vg�B���n3���7۾�d�h�G�zW_�]�-i����/� ����\�e�bD& �MY�H٫&�F��^�c4�{�5�J���
H����JX�q�$�XL�F�ăhlIh�ꭽ���h�w�c�|�F����E1�n�W�IVI���r�<�����Չ�kz�g���V7�/
�5�*�qU�>��,!Q�����^���Œ1�����`��Z(�V�1�b/AW®tp=W�������P�7���W��v�,�n`�����u,Z�)�j:Q- �����t*�z�y�no=Y���V��B�668J�J�{�@�������yrŷ�w_��8�y�°o�V:��;��ß�8<���Æ7OR�}a�"%G���)��_*��AUT����#���$
}o�uq��+U`��{�@]7\N�8�1� _$��"����OϿ���6%p�xG���A=w��}-/��a��}���[�>�n�I����c������tx���4*Am��K)����t�7�����P��I�?׭"R΁�`v��׬���鑴2���/��EDs��R�ոEF�.&#9l��\i?��2f��1�k[�>l|�w3�o(�+����uޤ�d�&>��P�e���I��+ݨ�2��~p-��Y�]�n��+�5"�bZS���^6���Bm�*��Z	Z��U%�k�r׵_k�:�=��=�C��T����f;_|��xӉ��q�v���ȃc#;�	�(1XP�6x
q����T����T4��4X3n倗��tq��p٠�0<'0(g)oF���07Q_,�.=�U�s��}�Q
�	��t%�Y�s�*W#FP`䏴ՙS�42=V���-{~ɴ8�k����B�iRVz��z�[Eb�A��A���:���=̽	Pv���#�|��F�4b%��m��Z']�_K\�y�`D{|h�?�(�A�p�¾����J(����U�וe�hZ��nĳrsIo�7ls�ڂo�0�$��)�ڐz�E=�����WBYmA7�]�YRH��R^��C	��
p0�FEF���]`}������k��[j9��W��(󤫛�}��ckxK.z:��:�����@�z�Y�c+����sP���?�~�F��oP�{�wO>CD�<@:��#/��e�Ǵ>{^�u��A�H�R� �����0� o) ���,�FF>��:���0�K���5�}�.���s熟��-j��&m
��G �|����<|�;?޿���H�Ǭ~�����=�������䖆{���w�O;^|��A�+x���kdJ77mH���?=&<�m[��Iى�fl���&c�1��1�N���"�+ox����ɡkTVT`TL9�1�;���?;�ri5�ˋ����ֻ �_���3�o��ǳY�q'� $/ꞱQ�� Qj�uv�F� Mq����*5�5sՌq��c�� ��"���hSކB�Zc\b��y�M�3�Fo�(��騇������
�P]Ft�A��!:�Nb@��0���Q����+�����;�-�v�n��D&�b���c��x�7C|A�8&_�+�w��Cw-��߰�ְ�>�Da�k��_����4P_Uy����پ�+B�oZ�����^���Li��Lo�����,)Q���5b�'"7��E�卶r��br�_^_�����`.�!�S��9"Fc7���q�xЩ[̚:+���~��>��Z�B(��p�{`���b�]�eQ�ps����7�0OSB����S�mPJ�0su�*v-�n~�o�^NS sh"V�����r���{�̬��u��� X��skzkB�E.?`x���t+h�ս�
�l6�OE_���"�"�ۜ& -B�Q�[�Hoī=��Y��}��n�(y��7m�3����xi[���<���e����O�1?�Gw3�����Z�|h����.���Ru��H���X ?���K#�5!9м{{A�O�5�U��_���8����u�S���L8X�vmx���C�������ej�	0�a���?����6P�/Ѧu�?.�6���\�"s�l�P���Њ�6C}���č�6�g	�������3���-��F.HJ�m���0��1�.F�9H6�$�qb�R�i%�rM�#��՚�
&�chi^>��'�o|����֤o�y���i>��/�)8;�ɀ��P*x���۸k�(@r����ֱ�6m�B�:NK�-�=�qK"T
�x�}�y�zkͰ� r�}��>|�{�#K� �H�댏�.�{J�����Z7��
�%OAH��7��4�Ka��]�F��89^�	�3u ��7;��*�����t�6c��~�Ţ��;*_L�I�k?t+;D�+�4		Us���m0�h)m��&�`�J�d>8����������jAJE�`i�(j�O�)�N"�H���QĒ��{�7I�#(8�)�fd�as��%��TZ�����d&z�r�#������NOɵ:w��|2�Ӹ�Us��>�{����WW{��O��L�И�p�g"7ȡ��|Y�|�?�(�����w�^"jջ�/緹��[ُu5����ݤW4�PS�<�G4k:�Cڦ�=�Z�������
ǜ3j����\�.μ��)�%�)��P��(a��H7k�r��ꑚ;�L��c4De�ɱ)��y6E��|�k6�(�M�ӕ�L�	*��5�?��φ�|���w�X�tk�p+�q�\�o�{.�BnY�eYS�WDK�D������M �I�Ys=A�BW_+p� Ebz]9�-�f���Ǜ�J������Gh��5J�"��-j�W(��K�O~��c�.��[�(6����O=>��Ɖ�,�>�����̟��O鋾}x�����)5���Jr�Ǉ�jr� t��Y�7����	P��'{;�B��Ĺ���>�ܳe�����C�+��0�<vt8~��a���^hi�E�zvM��0L�p����*ty-�ZE*�Z����a��-D6q����箜N�x{�|��a0�-���D��wu��ؽ�S�ڷ��),q:Hv`c��Xi܆11{U�^(n��
/ 0=��ᦜ�k�M'O�L8W�R?}�T�M���|����Qڮ�"g�x���?�I¿<� ��s���pp�sϽ�0�QR�wD�믿��nݺ5���h�����p׍�k�-�U^�7kY3�{DN�g����O^���T��Y'��������"�Y�� �hr!	�+7�\���HY�8?��ui,�=����x�T�Ƅ�[E��v[��M
%
���,�&�j�c���\����Z�m��d��;!��u�[sN�������v��s=�o���r9�F����>����Ez�;f��I��m���3��Q
���|�H���,�&��̳��k륈*�X��QE�A���&˛��訁�5�o�x,�ֳǩ�#[Z����@��D��l)甴�+�yچݕw��&�=J�" �P��®m�{�N�مO�x����:
$Ta6�iE<ե���+KL����
�1��S'aJ{B��@����!��ߦVy�ҩ�F���ѐ�������oa��ڼ�w<��m�D��eYz���+�tF�ڔ��x�.02R��x�O�����&�G��Y����EǾx��o���J6��Ǐ'�y;���ԑ�0����dmMM6".�;��WQ
;BV��<>|鳟`�@��]B��޻cx�8�;ߝ���mU7��^�u�R����������D�.s=�9���Y�k����3?�i���=�P�׸S�����u=/��Y�H#fC�����g�n�Y_}��ч�J�s�>.�՞=}�����X�>��0	(K�ۀ CzR	��^	Zy�6�֡����8�d���]�az3�t�Wٛz�-�j��������E'q�w_�;��RN�V�c��2��u�.�s�N��e<�t��[W�
���n��C䣑,�׈R�������th$��)�s��w����5Ǣ����n�d�k�l@�[����u/�YN�c���4~3d�|�HP�5.sa�,ƹ8�>k]<	 ��q)��7O���NP`�]=ٙ��ФB�M;.Q_,1��;�b.|�9?A���E�u׉�ۗ�"or+_-�#"
����7�y���m5�E�y�R�	�s}�ō:Ǣ7���������)�ߌ������b�{u�yO���f[�G�G�"-�̄�*�R�]��?����-�PqLJ�E����b�sk�6�w�m�,��!G��hf@��E�x��He����;�vi�֕z��=G��5�ۯ�[�]��r�CzG���a{ CQ%ږ��Q��Lo�7���K����X�1�l3��%0v	$���[ J9t�p��֣L�ʑ���OT@a��nº��Z�56�w6�f��κ	n�v���@�V��!�P��[rd�:щ2F�'ᮢ������w߻��Z��G��v#H�3����G�G!��Ƌ�H��g��0Ϟ� �qc(�O|�I��_�X>9���?�yܲ}3����ȁ�a��㞓���4�x�����&�������{�� ~/�~�\�|��utػ�� �u\�E:D]&Up2i4���WV���R���\��7�.�����v@ͻ�Qy�'1�0��>gc!C�*o@�!�HJ�K���>�������d
L�������7m��22�,
}�*VE �U��M	(ح��*^��h�}MaV�qC�O<N��S�վ\�ߋ�+u�`|��ƙ���>�����;�9k������a������~�ϩ�ϝ;/^%�7B��o�K�����k�Nq�`bTX#Fzɯ
�&K:um셖W~X+}�y�?¸��`r�(�h=�uܖz�*6Z��rH4,��hY��)��')#[G�xU��O(����4�m�j�lU�d�w@/����xOw��b����u�8e#�F<����\~�Y��^��R�e�{���:_��r\?�f�7���@7�˾�~P���b�5���<��&�1E�%F�-Ѣy҇F��N~~�(t��A�����C�`o�23�_)��������-?�-�t:`�OdϗE6�A�BUڝ9�+��~o7���X�t����[�\�fh��.��j�����G<u�Ӆ[`Q����Y�e�S롗�\��uޢ���cu���R��R3�M��X�����*����ϧ����3�����n�ӛPN*_r�7�H'�/me��3wo�ܚQ���ث"���|<����]E*T�=ק������X�Ȉ�9k�y���G?�E��c�ޖ������5��o|�f-W��	?h���O<pװ�<�>j�=������H�����?HJ`#B�����	Ť�FB̀t4��[]�rz�z��p���BV�-_���	�TLw�&�?	�����j�f1n��矘Vi ��^�0!Wю	<�� �륺E`	��)��P�\���(����]����"`@�W`�KȚs^����>7��?�ï�G�,v�����l
������k�,4�[�(�+b#%l�W��j9ZX!N�x��jM�h��o��/�˽���z<�*����D>����Hw��um�u�}���������<J��~뷆�{��5���=�\�̿�G�1u�Y;eT9^�D7N>�[h�Q�牆Q��׈�l"Jt��=7���`+��HMzz�&%ʙ�����^ެ�짢�6���\��S>_sQ?��R������
sת)'c$"�h�^�~�sJ�Ǹ���_���Q�5e��i9������`oND��k=W��{.>��J���%�<��C:��l�Į���Y��O#���1��"w�BG�����K��e�,�n�L�h�Η����N9�A����hH��7y�7�z<�B����⡶ܕ�7���zۅ�A@?_)��L��(�����{��|�Ub���J�F[s�6�\�޽{�ε��9(�N�2�GE�G�ExՄ�IU�Q����O�a�!�^��׭ �Q"�c4���h�U[�҈}�r��hQ��]�|Kr���n��j��X���P(�Z�ʖ�©zo��?IL�f3���ն��ݸe����?�~��p��{���vv�P��Aj���u�	�k�b��رe��8m��:���Ƭ�׳J>Snup�[�D`vflطs˰o�f������O%�`��+���a��)��
�NB�I�����@t@�#�m�r0�bL_d� B=|�
�4�m\�ᚖ���5ap�5||��}ۇ9ش�	�?��/�0�{�]�wP���p����UfZ�Mo�l��1�!����o�*8�C�Ғ��ٸ=�n���es�0r��b��5o2
Y��t�o��o���
炈�n�t�rޖ͙G7'���`���o��o�*ٵ���?�����?�T�a~=��Q0:0���[��%T�;����[��U �*���v(c:���%�l��:t0-|Oѫ�ƕ����$�U��dHV�.���&{]㹸�E��{"�R�떉h�����1�k��g\h�)�M��7W���9+�E�O��<R�˿Tx�^_�)c�>��wߥ��,�Q��-]�ܑ�^@l�܂����¹T�K�Vi��{�E��ږ��MD�<�x���8r�k�q'>�c:��Bbw��)������n�(,חs3��Qd���@�6!��(�f�^���	�7?� 5��\�:���u�fH�FF7��*�\�n�[��d� l�Xs�������������C�>	���m�;�+�*���Ϝ�w�guғ�vh�T
���~���'A�ޤ�ZZ��Dy߲Fk�l�[xL�+�&���8����ǌ���� ��:V(��,���Av^��f��{�}��-�#J��-��*��E���ί�Xfvf?Cx{nx��w��(�x��C4��v� �
����1_�{�-+�w��&*s�#`��K���]��jt��� �e
C��m�Ƕ��nڻ~�Ệ};T���/P����7��4���)_�F���(X��߂���D1�W���q|�!bDJ�_&��2O�h�Gț������͖?��<�;��&"�v;�A�s�P�����l���l���VCv��102�����4
�̈��s_ۣ�tv6�{�n�s��\� @��5�mKW���p(%��8M�َk�4��w�}�N���[���{�{«�?
�Ν;#+zw8C�K���.�F�Y��?���i,}0��(^ߟ=��>
(�s�1�F�~��50T����A������ʐ���"/·�S��(c���Y��g��M��ɦu�T�>�3�7���,�ri^w*���_��x�m�� *bX��jV5Wt_�۔��ټ�;4����=(��d<�eqe�z]��G�s��_E���˟�RZ�c��M��P��j�@��k���+�j<��C����Z�����(�UWmu�nҮ�no
��z�j�`S�0����o�Q��?������=?߅A���[�Џ;*$Fa?F7t��)4քb	I��
�E��+]"�4���l�?�Nݻc�p�&%�+�l����T��p��p���6Qص}�p� yG6�['N��C#�'�v��ݥid�5�= �>K�Q;��Ү�iK���3�"n�f��m⡇ڻ���Y�	��Q,�9E���H
�����?����fw�!�p}8rx�p�й�����I�[��u<C��i��ѷ	S_B�V7�!���Z�	[5� �	�z߈
��K�9�V�o-O�s`����y�Y�֍�$>S(���w�������h�s�:Áh�ٍJ�gO=;����*�-n���]KNr{~8�o�h�V)����R���hN�q;Ƚ�o��<h#�P^�B5C[�M ����nb45�Ԓ�7H��A�T��9�Q���}�����]�T�ɏ�Z��5:�#���jѺ����U�7h���p��)�	|=��6�ƹ��5Q�ʖ.�R��?y������G��tע�9j�e�uv��0j�����Q��R�DalK@��t������������.>�{�	�d�e��l���c�(?J;K��Yq�s ^���2�Q���V�S��R§-1*ڢ-����P��{��Q���ɾ̚)o=�ʳ22Jn�����7�F>;5yss�`}֑4NZ$4��KK��~�:��FD����M5�e�o��T	P�:��:���Awd��Nnl�P[J�>(����f��bM�M�׶�*���2эW�j�u�}5��2J�t��c�V3 |>z]=?���2����qG��hnԋ��O������W���%D���
�`������,ex��������J���ײ�������˿���w~���� l2=��~{��o=�]���KU8��Q��Vm��Sl"Ѹ�2���u�g��R�+�2�e�!lJ$�$}Y�e�7��&2j]��O�y��̰�u�R�g^<6������ �]'�2���a���U�<l#��H�۳-�����7#`,����\C��S�fl���5���MYP�w�OOu���Mݲ�ĺ�nnӖ���
���;��T��47L��4|����7�7�^�N?:��ҋ��I`��q�,:���j�eв���MflU�����O~�>��)�C�.���#�:Rh�_>���s����Q��_��Gk/vƶ5�u��{4rE��NCjd(մA�����d4�N�@�����U������|���'w�a�
�P{7��LH9*�ei��h��}ͰY��O9��%� jE�a�8���=4$� S��S�yLgC޳\O<O��k}���>c?a�1*T���S�ҫ=��R��3|:֞K�����q�K�b��V$A���K��h��8$�d�ƃ����g���Ջ�,2^��@DO��i
��Ƚ��R��d���ߺ��z��0Y��qݻ/m���w��_���;��W)��_����C���L�R�n�[�]Q�z��F��׭ U���J_�i7\�!�������������z��������]P�U!�l��F=�n��ޛ�x�_�����֊h�f����7���~�f&o�?�c�y-�pѐ-�mt�?�����������~틠�g��{�G�Y��K��rnzۅl����zЅ���0�n�Ox�����"5TQ؊��n	�dZ[}V��۱j�Z���;Ǉ�����S�%�?��q������B/G�F�eI�U��%� ��s~��ru���DX�&�]�(��0Sy�#��m��=ÉS硚}���	�n�p��$��Mx�� eYi]���ؘ����ר�>2|ꓟv��7��޻��edx-���]x�@�Mn�h��ER"0��ّm��i<�bP�%|�s��\�
�����Djv��5|�����/��] �9�� �u�q�GgyT�}�;U�s{29��k�㬳.���`8�!�3\Iʱn5jԍ����L�ݣG�����T�e�B[�6���~�%�Ͼ՛cz�/[�4O�����p��<��0���v�}o�W4|������0o�1�u�U�ݵl��q��y܃g��Z�Y������:|	x��c���V�o��&T��S�T��Ζ�aٮ�ͫ0�t��7��=g՘e~,]c���2p�|��j��viʚ�&8���2��`+�:��o8�(\��/�<ɽQ����i;;��v�Yw��W�{*X�`�}1@[YH�K�z�,�K���[E�D6�aKl/�7�Ք��z�j��D��|���FI�T.#�&'�n2oW�����
<�+}�����66��h����G�ص!��e�<i�[ϑu��n���\{x������u�н�Qo9ۢy>�!����u�r4��?߿�?3������y,�;���>:< %�|��ָ��7!��I��Y��4�_��}cQ+�(�ϧ��A��A������g��9rǗL�aL37E�^gдQ��Jd�t��x[n{�h�Bj��#X�Ӷ��筀!�܎������/\{�rϗ�^@#��]���G}����3x��gO��6d=9��1�vQ��q�x* .]�Fkǭ4����>���G���0 �zr���_��_�{�[���l��ȯ�n}�|������5v���/V.#�P�x��	��^v/�)*�)��~�4��8�,\ ��ֽ���wx�����Fʤ7�x	e!�(z5�Rd"�-{��-����������`�_g�N�-0��ݲ�~LĲ���!�[�W��<�����YC�b2�77��R��&J$X�2���Ͼg�am:]7���={�D�-A'|��6JU�7��{s�/��O~�c<����U����Z�����h�L���{��dS�9��FJ�D�[�nOo�/�6��r*[\g(m���c�ZY���!�j!�!S�1�A �Mz!\��L4a� ����.���>֣t�`���q��8�[�}�S�(�µ�b�����W���0�;%�ڸ�fƎ%о��{>y���{��'�
�b��$B#Xͮj��=�W�N��p2��T�{D'}��g�y^)��}L�J0j�Q�u�C�lE�-n�*��s�Z(�K#V`�b�/I��O�$`\��K81���nxY����e���W�%�u}G(tۦ�����)i(�`X�G�3d���p��mH�q#�k�)��q-��J��(b�U�������!�
�U\�{��~��*Pםm�wME�4�+��Χ�{�l4"0���itO��u�~?�u�
y�g��� �����4j��};�6kmA_o$7ڕg��k1�/�?��	�mg�Y�0�-<�}j|K�Wc�r��k�f-��u衏�ٞ��Q-�^��R.����̡�b�\}B+k�}��gs'���_p�J~Ae�W�P��Ye4~�^J����C�!���}N�7���� l*���ܗ�����-�6�x�
����ϜZ�z�9x�Y��?��? Ran�B�Ρ��x������K/��f	O��h�������3燧�r��q�|v�ҳI�#Nuy��I;�N�7}��(=t�$����~�l����r� �T��������0�M&�z��^"Mq�:w��BC�Ϟk7H����W]ʲB1T���	o��.���7��K/z~~nx���
{۶�	���1�~5��~����)s٘��U�~�*ts�c�4��E�\�.�B_�1�s������J���eª��F�Ч�;ʯ[�GTN����P�>������˯�!��ڸ��&���	/���L�A�u�^5�S�1S"��+G��[�i�Ҕ��<v6I�t��������c�����Ki�깍�X��PІ���(t�m�l�����95�7p�(e��C0C�IbR�s�wf�C����vu�u&#�^�F��Zf�<��g�o९g�\.3f�Sx�IePwʫ��
�
<�����9~���ϟߨ��W)�:�5�����ە�h.�a}�?�P�h���g�
�!��P>k;��Yx�y�	�y"�JД ����Q�|�����Vs~�/��[YJ�H4zz�$��$f1̥�+�3��Ր���n����.��n۾u�qe���Lʦ�)�m�"�6�%��%��"�eU�G��_�R�.4�35�\�p3筷" ���3�
���}��/������o�XZێ}��׋�d�#�!
>���.<�i`�1�۟ky�8�xN�t��7��<��ؐǈx��L�2�L�����U�����+�Ϝ{�p�L�4�
${���\�vO�R�#=����÷����ЃSQd��W�-�ҵE�f��\�K 	�- )>���&A-"#�8��+ MF��\��@�� fn��	x���o�8;��{�~�Y�^ZAK�ת�|�y�-��x�`=e\���Py�Z�G�X"(F��[��]�"���{4*�\��[�p�H�ji�� �����0���zr����o{I"���/�"�z��1 F���{�ˈ9���fa�#���:���>j�/�e^r��ި��� S�f]C��a_u����7��ؓT�\�L�����:�'��� �Z�U΁�[G�r��|U Ďu�TY+�3U��s����cgiժw��hߖS�G҂��F?���-Nf�m`G�Kl���<N�b�A��9��t׺ڻ�tuH�0<�o��P��x6*bT�e��F@����i~��կ�Ɨ�O��S`}ڍ��w�9� Cy4¨H�6.cD�n�4RH4��'Bb�"�X�������kyF]������:g�'���M-� "W��kn�
�S��H��g�w䆫�N)뎦�������9�������tEdv)�B��
ܩE�r)~�gz�����[5� �'B�m��=7���ٗ�W���|��# �����h���$U�;���c��8�Y�Gp�q?�!j�F��"F�X��n����-� ��Ƚ%�g�K��X	���E���6kg����S�4%�ؑG^���N/�OaE�M�VC�K��ϡlqu�Z!��,
\����4�Y���5�w�|���뷇̈́z�Onx ��ÃG?��χ��.��we��{_��'���C����e^�c�Bs��q��<�Y�C��Q%f8���&Ü+�k��p���$��s�
��̪���5�m����Fhĺ����FV��S��UE&�󺥝���Z�Q�%�/Ɣ���\r���4���6"J{U���1b�=��=�M[*Iic�y�2�z�E�\���ź��H?��b>�A��^�ىiV�U�K�m8����#G���q���s�o�k��~�����);���� ���AJwV`�MZ����1p?��G�@gv#@8A_l������@E��-�@�#b�ޔ�:+ݬ�D۲t�����{8���$R���/%��������n8�u:+J�s�Ȝ���r�*��0 p2�eK_�A�ԛ�"��DO\���s���%�$g2u���Έ�ն8�~��ᕗ^.\<Gl��я�����9�{y��+�n!@f>eD,?�#��A��PC����x�:��>�;Fi�y�,��iQx�uZ+)�BGi���&,�x�=��Ӈ�o����[�a����5�[m�(�4�(��[��t/�pV	ʘ~��F" �e�5���g~�_�j��ЮA���m�K�ݕ7%p��z_��X��{/Jo'!M�va�i�B���h��W��f�d���
�*�� �s�P�5끱�R>R@!ˢ�VƉ�R��z���������1>ڕ��X�e�!AS���>�я �"׆!���/j#���u�� ��x���ُ>B,<�y��:Ы[��	ᎍBlbry8t׮᭷^O>w�P�ۇ�ss���9̢h�y���"�˒�,"X��?@�pWB��6�nϽ���U_{�V���r꺩B�u�R��88o奲��b�s�r5*`O���4� ���jc�w�][�s�<���Lx梢XkzA漛Kx^(��2iq*𫕒i����(�n
��"�[��*�[��]!�G��M[�q\]�=�$��6ڞHڠ�ٟ�Ǽ�N �T9�� _Ŝ8$����a��k1*/{$��w��.��[5�c,U4n��&��c���Ű9���b���H�l�Yˆ�3�w��1�sx���a����ṗ_.B�,�KQQ����h�u���������2����pP�e��[���#��]�"E,
r�����3��.^=���f�y�sMkh] �r	�}9�O�:�{�N4`�u`EMR��e���s	�s��ft�"N�k�6���d��w��sx�q����k��Q���X C�n���އy�%�o9�Ir+����" J�s�$���#��#��s6֮��>��? ț ��Qm�+�nߊ����mu�eE�T�������2�f'kg���s�)��ZM�T{�s=�f����f��hRX9���w�C/�G�lZ]l_���`�z��)���]��N�"̇Ww��S�}�P��m8�Ojbϱ)i\!��_i��uz$��m�w�Ǻ�j_� ��|Z���Sc�T��<�֌"�o�aT`¹*C,�临s�2T�;9~�A�y��(���T��76�g�n����<;<	����=4D�~d?�����˶m;#��1_����������7�7���ςt�}��hn��j��n�lټ�\9�0xЏ?~������6�˞@���`��W�ܕ2�J�Nzz']�ҧ�J,�r��kߑq��Z�QGO $�)�Є⽄���4ү<���j�-�g��|`��S�	��.n�ǐmt=KD����mD2����������2�cIQz4�\�%��'/\Q��T?O��O��ؕc�p���MŰm��TYx�}Ҵ�����/�@�6�`�Ɯ�4�*c1'��� �^P�*}���R|�׹�{w����~ޭ��HKk�RX������z�}��5xMFcV?��3�e�]!�}��9s������!R7FgX��bd�}����P����#=�Q�PK�V�T帷���I�"j�G���������0�)��m�bӤ�Rk������笖G�B�e1��+�רܸ|�"J�<ǆ����({@��V�H*�5���U�P,eX j��Y���,��")�i�?�#�����"7xq+�RX6:�����Snq?D��%��kb�Zl��N�uG(�3g�<�BO���+�����z�iS��6⡛�r+&�Y��*�X��+���9�icu!��fߕ�6��c���s���Lj#զ�{���;�4��{�B�!�<��z��Mx�?J3���B���`���Xʆ�@�^Z��� ��g7lb���>	��1Pۻ��n�]-����t�76�̆1:�m�x�}V�8%<����j��eNeP��7� ��5�F7�F��品)��Q݋��Nݓ�ס@�GP?���^Ν;3�w�����'N�&���]Ò�I�Ɵ}����[��O�n���$�~�zB����p��"����'��>|/��pE�;}�8��ΟG��$��j��'������������"�ERQZ��Ly��1�w*ʤ'cX���
zh�y^��}��s2��642.
�r������n��H�R�Q�#�L  ׬�_On}3�Ķm;�Ӕ�A�*P�9ī#^ߖWh���:sN���(`�����|��.i��uDy!�ס�r�
��`���a��O�� ���} �>ɹn���3�=֌Q�������W^ɱ��և�MYT�2��L�YI���=��B�Y��+�h�NX-Ӎ��ze���.v�,��9���,l-w������NA&$���mɟ�h*��>����6��������SI�ŕ�
['"�ܽS2$��Wբ2Ճ�ܠ7�R��:a�ײ4s~�,�n��>�T��l��c��2�������w�?���`"(�q��u��
Q�MD��Ll�>���?}���J"u��@���J�	4���A�,�X��LDjy��Z|�9� ;��&;R7��R�"���
�f,��_�˻��|U��M�W��G|���"��;Z�Z�Z��_�Th���Clk��&t�'\@���� "@ݿ�6��iJJ�VK�l9MYp�������[��ZN��H�.��������^}�J	��sӊp�w��Ʊ�o_%4��{�j|���sj8v�,�׭��]0�ɾ�&�j-��]z`�|�:���p��C!����r���gtUEZ!��t@�E!��ߚ�^5�F���Uom��ֆ��`UI2V�Q΄w��a�޻�m�ۆ?����e��D��$>t� ���{|����\,��#�5���mG�T�voR�2S9**s�zW��%���T�m���9"�����3���֕F��X��EB��[��x�έ�h/�r.}�υ�Ӛer�1gT���w�x�25N��c���i�#+[^���3ˏT 7m8�o�q�hog=�{�ܮ�q7�*���LM�[e�rDs�^\v���Q���C��*�E��8[ޫƶ�c�N�I��(�E�]o[e�O��=�r(t{֠;F}�o9�=��g?[�|�zT�6e�����!�M��j��e^�zu��!2���Ip�U��~�a���I�b��2I�<��"(|���x�W�ȉ�B����4�=},J�,�5���ƧX�V���$� ��S�Q�� �Z��i��0R!�q����
���-��#wz*����T���62�<�D5cD�1;IYޖ����w�� w�p���ͷ���b����ڹ;�����4.+��!geEpB�Ş���T2��NX�Ls�� �R����H9.r���k���<P�S�3ރ Ks��J@�EZ�s�W���\�!�p�v�U�����T��S��p�:�E)X��	���������?�R�ցy�]q��v/~.LX-�չ��ZW1'�Y�OO�ŞZ���.G=��Ʃ�o�p�I-ߚGIlH�j�Q�P�r�����OH��
���m�=KxT�Q$2�ݦ��p���]�B��j�8B�{HZ��RA/}\����\�%4���!�Ǫ��{+߷�ښѓ�ݷ�9Of�a��C�G��|�r������e��SAn_��֕݋x	�	��MO�p߹D'�˷��4O�>B������w�'�Ͻ'���V���5t�|T
ȉ25�D)oU��"ԩ5|e�c�f�_�����.�w�����w�Ee 9jR�_�.zzZ�=�6󻛶�2�۶��Hv�|�k7�����w���
k#T�՛ẁ�Q1w�������?�P���u �RV�[���M�Q�_�җ��=?����~Ơ�4�/�9����>|�p�ǽ����tf;x�`�D�خ�͛[�.�1<�q�FdMS��=�X**rRh}��B�:�A�Q�������	�)�8K>)�Ҡ�-�-�#�|�=*Q�'Ξ��Q� Ϊ¡yԆ֙v#oF�R�b/��G�?E��<)�E��b�~���ĳ s�DU�H�sF2�m�3��2zȻ��dcM{)���~���(w90h^�yv���C�'N�����~�I6��(H�(�m�Ml�_
�N����)���%ݓh�t�|���d6��	@��k�~Y�Ub�s���{�֠�����]X����M��4d��js����J���>���-g���u^�|���Ek{�cv
��q6���Z���%\`Z˱��܅�����GN�*�	���b���Q�w�y+��'��cTN�SNzIn��`�?/�{7��� �*�����ق�ۏ�|=J`7V��,K����+g�#�n��y��"��*��P�lS�b��5���ꡊM���/��z8׹�z�l�h�.+x��H�iSr�0=z���g?�	�k�W��5�x��g�W�=?� t�G��ko�z��p���{�`k����t�b����x�g�_z�<��tM�Rr4C�6y�n�jX�s���6�R��������E}Ҕz�K�oW��QЈM;��s�Ʃ�1k�v�X��2���:��N�J	�]�S.��u>���}���Í �(9�[O�\�PS �����Q�=e��K��<���<W�T���1 O�	B�c�NA �kV��P��+�����%j���y�Uu�4?A��iM��H�ֽ˦<��?��ᩧ��5\�ç>���պA�z!���hL�^^�u�΅����a����^KeI�,�3�l�����N���9�V��S��%4Gj̞ ���l.�����������s��"SOz���sou�խ�4~���';����3,ş�531��͉�S!�l{?�:�G����4JR'Kz�Bn%�������)Р���|2\�0g��L�X�
嬍Y:�>���wh��j�@�9
ގ�\�ԯ�������3_���Q���L�y�kJv��tp�K���7��%]����Q����2����1�k�rh=̷F@SԅO�jJ��(j�`?�r��s�uW�w��\q]W�C���̾���&�^��l��ּ�|�+Jx��a�u*�q�P��7<{�w��ل��|d����?�DاކDe^�V��%������/㼜<���l��cg����.�R�J�"�f����@�������.��rk��5���RM(s#@:��gl&�2?�2�ַ~2��HD��������>w�(E�ɻ����S�����a�7�z�?x�p`��E9\%���5�	#����s����mÏir�}a~p(tǡ�=z��p�<@'�����H�2�����DzJ�V����?uo}���+�[�~M��sX��G)FaS6��1�Z2�Ud#�'���[�����Uۇ	������a<���!��#��5��ZR��/���`ޗ�(u����hz���l�F�D��D9��Vqv,L�Q��7����}��P��ӷ��}�N�{=�֍��Y��Z7J���~4�ѽ��.���2�O/k���p���|yf3�݁~�z[N�oi��@b(��jD�d2dD2�m���G0'gUWA���V��-E�<Y���JmY9!�����U�1J1�E�}e�16*���f �����LJ���X�_|��U�֣�+��\UfDC�� M]W��?�U2�j�Ү��q�05YkVT�ڒ��r�D)��"2�1q̲8�kʥ�C
����%���1" �_~u�:s�{k���4���Rv���x{�΍����B1��{μ�����Bq5�ߔa?��@��m�c���7a�l�2`�r�.�)��'�7?eN� ��eyf�g����-Q[���e\ʡ{�i��Z�Bp�!@��\si���;Gy�g���������3}���w�����?����g�C�JJr3�M�lm�I)'�����o��mO�|�������αТ����FěWQGn� ^ۘ%l�l¯{D}�z�aU�	����|;f̬��lt��E>���ڸ�p��~�0A[��k7�M��ax 2Y|��q�����;H�ov�����(��D*���P�|�^��%�!������a�{�O�3��#��y�ҕ��#`�� ������M���C��t*]�z�5�N)�R�k���|�s�:C�d�B�ѕj���gZ�b�lhpp�S �'	�&="�&�=�z�!;�ځO��2(rrג
͐�zz����i5)3��l���Rr�%��='ajäajc�̑�z�5C��My�֋w������W� ��a��n��+��݇rè]�&-`w<��xe����R-"�>K�u}�G����&L�x~��Mi�B	I����Y�&�{ɩpP�7q.I9��Xq2����3i����8��FA��|��� ʕ����6\�Y�ab�=�r�4�̌M�4o���Zn�Βk����S��=���P��X���
4Jf ����Mos�+�{����>M����|hЅ�^
�nql��`��0�}�m�tם�l�,��$ę���'�vX]���o�B��c`�MZ��������/S�<�R����J�B�6r卺�ݰNg��G��g���͔������&A7á�[9�`�����л���aʛ�`p3&Z���T_{��J�Ɖ�w�6M/�®�:W'�螺���Z
���w�4c��P����_�����������=>|�?�\dr؎�����j	��畅��̮�����aw�:�����Q
��Q�S�Ү=����5OsT��6��hj�CeT�y��U,�\=�Z+FSd�ByM"<�Pq��e�wx��O�tt�D�r�z�1�x��i��w���"B�'?{a�v�2�y�>x�o���#�w����e��+����|�QhUOsN���<��ZO��}D�����T_Ö%�Ǩ�^स-YJ՛y�<b�A__�%��fx緓"���K-��#���	�p��В���Si�{^��4+��y�*k�G��ʡ���1��쑶=���(��U�A�Ⱦ���s��#�9Rk��!�,���wc�˓��F���B�G�=�vT��T������'(���xW��37�!;�C���b�B��?�1�/~k��_���p�VV�+��m�R��:�*W/��]阤ɍ��5�������FZ#@2�+�A�e8�H78��
Y��5ra���o���Qn��D�lq�8����F�d���H������4�����9m�i�|r�e~OM�&�1�4��9ڬ�f^���0�:=9}}���DP~exܝ���
e>��:!�C�yB�YL�lkU#�_�X.��̟�O��B�k�. ���7��A[�ϒ~=t7z�\����~U}v1m����ũ�f��"J=�t��P�
��W��r�����x/��&XFQ�U�ܬ!~Yb�P[��區��|s��?q�������+Ã�߃��cSA*�y���G��Ͼ���ir�z2vW��(�'�9�#_�|����kx�����}�P�lKK��tn��ix�]�����G�B�Ѧ�� ��Yb�MJ�e�s�?Ԗ͛�d�w�����A�� H��x�s���_��_����Q��>�7Ets�"���ӝ��Y�ǆ��憓��"�0v8�5���Lo;b��A���|fEՍ����u��o4\���w[Qh#z�q�أj}mEV��0#5n~�~�)+���D��>�:_?W�f�W1���s�����Q��ڃ�Ǩ��s5e\�R�JԆ{L�Q~w�܍�j������xu�=A��``��J>���*`���.8�{2J�Bc�K4�Y�N_��
�<�x��u��*����Q����\���$��k*��eO,�[��0��<�g)��~��P=	L��d��r���.�yE�:t'�����a��&92���&�����+
ԁ���/1?�5��SsD���O���C��Y��>�(�]>�k ����=`�1X0S$".��O�y��*+34x
�D����إ�2cB-�T֍��+�:5��6���y,*:�Oڕ��W�K�B/^�*�"Y����	��ԡ6y����jFC����\3&�<���,%t��6r���Wy�������ǝ�SǪ�e�{�J)���+d֭i�k���6�߽:/,��D5�p,�1�h�в�G} ����
ݟ �	�:t��a��Y��o�V��h4�%o���������α������^ĳ�D��B�(:�����w���|h�tZ�>�m����{,��ͨ��4�J���LِR0�~�k�~;y�4΀|�N��������ʅ��RΡ��"�,��kO�v�5�H�iD;l�=��sk��m�<u�*y�R������6K���z���Rxױ��ڐD�`1�T�� U�5�1��)���T�.LyFx��(�}��#����"�%V�@��:��.�hĪ<슆%E�wM��>�����hV)�5,@E�T�������wϹ{�l&���D���kc�#{�{�m
3�>�a5kꑀ(�6c)!m�be�+��5KT뽢�'���-O�I�����>�;~���ʔ�a]z{��M)\�5��	'��x�z���`��yd����j2F٤�d*3s\Q��COz=�����b��{����s5��<s}������*״]�i��9�U�)sl�<�/]Μ� ���p�'Z2V:�#+E6��+e'@�h���z��8��}��Np4�Q�Sj{���9��^��˝���x�n��iEq�t�*I���Vo�O˥��9e@n|>iɚ���R������*���??�������y'e)�.��F$k)�ch�f	��{k�i	l_QTA '�)y����%)�>���zt�����P
b��
\����b�,ky����Ob�9��ޠ��n�P�`�+;}�t��NQʶ�4�y��%�X3��07"�� �>j8F�>D��=F*`�UJ��=�]Uޣ�է�r轼�MY��T<	W�sm��n I��6֓yS�Ҩ�UFEnb���ю�.ӣٶ�-L��z:��h^B����*%��=�F���t�����Ի��^m�_OuYԾߌ��F#k�"Z.�>>�H`�%Kr�w�Do�K�(��<���h���HS��Q�az|�h��K0�k�w�olM��e�c�T���b�O��t�X�{�Ae��Ux�GBۮ$�K�޶�✶�(�`�ۢ����ާ��{����!�ƷzZ�_�&!�Am�"����?��9����
�������Mb�t����hY����5���3g����F5�VQ)SqQmkժ	�JG��3:�	��Gj)_ݏ䶎�bo�1R����V]E�z0m�۞���H�^k4K�p�f���@�V�kx�ļ��M�7=&��Zr�L�\�``߀��=\�z����.ڤH����Fjh�T�����o�B�r��y�ڟ��i��.&�֖z�i|���bv;s��Y�-$������.8������~yM�Dh�Φh�7�p��>���)!ַI���ؾ[a�zV��UY��e����QF�E�W�~�1�u�q��b���1��w?����~E.��5���m�ַ�v.K�9�?NC��I�S@U[6A�I.+�AE�f#�E�P��@@��(3 z���5��:>#-��������f<y�2�����;k{oFa5χk�h����H0�P��@��WB�z�M�I��egT�el\�u��=�Tv�J�ܐ{u�?&��T 7��+���y[3��B�z�.�&l�zZ�Vk�4��¡|�cN
cQM^<τh`��1��5���m*m�6�I;;c~ݨԜ��6;��S
��H3>�;����^݃	�Σ{��*m+��P1���]%\��|u��XZ��?�Ԅ��	����)�B����	�O�������
�I�*���zծ�%<r��_#�B����^7��:��m<*���)'t�Z�Жr}�9��w��-��.��B�1� ��K��\L�u�q",R-��^q�'�@e�"_*_���a�X��,�+�a����^���WC�d�bn�P;�1oB�{��9N�H)��a�^��%d
�G�;M=9Y]v�>*�	]Y?�IOl05��b�!(}o��톗���Nw�A)�p!��۸@���L�R���
�Eu���ѣ�=��#�v�%�-K���^8�'�Sea*����j�Py5��l�2˴=��%dz(�^[n��[vUx&�[���E4���j0DpU�U���m(Y��R��$���u�Ⱥ�ٮJ�U=p]S�ڇÐu�Eh☨���_^���\d����,M*u�^�C�bG%�)��^}���|�M&$@�R`��{;J����	��̦�k��Μ;�/�yj�}P�NTh�<��S.����",9�"�Uw]���ސȩ6h^o�n���d�&8Q:�!�Lad����g���K8��)�*"o��pl��W�Q�"z5����A�./�6�h�7�h�ʻ���O�Ys?m�eR�km��(�����ϭ�mK[\��Y?͐qB^��ܯ�$*L<t�Ή�78�!�Y<F8��K��/�YI@��f��$��2�{>����;��<���nh���K����{��v?f���ki�"s_��<�2��x���9�EO������ն1����iH���R�#�5n? ��k���C�޽��s*��+Dk�����'��K0⥏���m]ז4���� (lFf��Pk�)*CNe�m�v*O ����3�z�<�7���j^Rk,K�-��e{���4P&�Ȼzm�tq�J���o/B�;sȆ9�k�g���9p���x�<QRx�a��]#���q��Q����iC|.�c�ųW���&�u5y��̉{LB"C�v���!��3�\�ק!��s���D)�hJ�����I�%,:J�I~���j����. ���޾}�y�Q^���WA^�-�x�ݹzoL�
OB�X�.Feg�^)6y�K��քf)��~rj��Z�Uy���V.�_��J���%�ʫi���T(
��!���C�B��6[)�R>�g7_��X��������F�<��M*��?;�ִd�)��˦��'�@�{MH��3�۶��{�ߤ>���,��T�7K_�^��u��
P6��@�Z�@v�R�ʏR��Gگݼ#�Z�PRy���ѨK�Om�* �c���lZ����W�s��{��a³�'#�6��&�<����Jr��~T����/��.���`��gT�/���}h�;�QcR�q��￴n��w�W��<f�Wj��J�����<�0ev��u����̺?4�g��)ˮ4�Q27�qZf��M�]e�����s2��v)L@�k���5����X��8 A���2�;kZ�r�
����F���c.o<���_5�뚺������fhTX�;}���r�+}��w}/�9~Vw[��zP��A!7��N�UqKh!k��׾�ȷ��&MaҔ�2FE�܆���Ŷ85�-�z�=����� �LЪ![����p���-�YO��fY�LJa���(ps�!���K7�ٴL;9�?q@�>�E���W��G��dm�����)�6���H[����d+��睂��7U�e��xV ����FoH���ۉ~�=���j!�]�:�؛/���E�_?v�'�U{����UٔZ6�ĄMF0�vSx��v��\t���_^y���th���U�>
P��l�'U&����y(Z�10*�ݏ��S�j�\��%j��m�z��Qǭ�o��n����cc4gY�uab	� ��A�ڰb�^Hb؀�傈.�c�M���CW������ȩ�7�S����=6?��z2���F;x��
��Bz��+]�ڍ���{ }"�Z�l�B);���S�4�����c͛�^A��B�"{�oC2��0��ǉg�G��q���4��R��L'V9�7\���*V �o�{R��/�~5=���z�i�#���[e�Ե��e��(���
r-z�2m�U�YEq�P�T�i�'W�{-|ֺk��5�Z�)c����r޺�j_<���j�3�BʵY#{;��Ws�μ\@n���`��x�Kq�5��汃$;m�,c=Џ�g�r��d���-K,�n����Q�F��+�ןj���^>L�;��W�n��[6��KM���	ʫnB�R���%�������҂��#���&3e��m�yx�Y*�m��s6b4y�%�4�z�\zO��et�,��7�~���;ÿ��?����ȅ����x"5��?��&A�Oo�gh�D��,q�݊r��30�M@_;�ޛ�^~�,kCp�DL��m�k��	��d����q�J�D��g�Ƙo�R�5Cwc�4��_nz	��"�^1߹�My�M�_em�J���>��+t/���CG?����>��G�6%X�E�4kcv[݄V����&�`r�Γ�
AB}#V��݁
�*p�KU��4)�ڿ�߫�s�.�VC�K�ӂ�X9b��{[S�=4�OX�#&ESh֌w�VB��R�ȚR�p*!���ߍQ��w���}���n�������y8|�a8��9�;A;���*���i6�`8��oË�lF�t�Nf ���)��<*��Q�y�yTR\��cZ7����v������3N�kc/��-��!��X'�ە��Ä$׳��P��'J�NP�FAX�[��Խ�&p[�fdI���S��mf�a���J�u���rƨw��F�:F��wM�B�R��R�ˆ��AY�/�/ ����V�š�5��~����s��(�j#�c���ɨ�l7�_�^�ųF��a�ʜ�~�O��z��$��:�F���q��t��^K��t55V��bX*��+�>U��y|O�6bX��wc��^�㔜{���cu�ܿ�e�����e�6D���X�\�+�*gL�AnkX= &!��>�1�-T�CC��`��K�?;���2�ub��*�uQ��x%�aD�h�/j����N��6�n?{k���M��Y�SP������o��_C�&O/=�S��<���;  � vk�7�%͞��nn�A�r�4w�n�ȟF�4��8��<�8������X�ʍU����w"�M��U#ZC�K�#{�{ǨY!2�����Fd��7��=��n�S_�#���;����?��z��=y��}e�ڮ0k���pvE��	@��(��5r6��<�EQH�� =B	=����Z݊��̇@6v��k�W����B���c�s���n���	�g����,WJ2��#^���4ή��M�F�.7�@aQo����5���ۄ��<m���_�:]������#�
|賳�C�)��B��nH<�T��f'����Z�BF/21����.�T��K�l^�jv���~j�k�x�M��C��i�;��7�:>���2��+�ʣ��Oמf(��Nb����$��Dq�[gw*�+�޽��t���HJ��+�c=��$��,�I�
j�����%�]�\��E2{�QT
"8�'[�YE��z��.e��d^�:�*�*���bj�� 3Ӎ���b�FU�v���2/]%Iŋ� ����K�����\�,��U�dH��hZS�}-�*G�"
��\�H׀��^�TT0����m�w�0G��j��?4fF�p{Wv݃U���y��2��L�w�^��52�'��S���q�0�:X�1�Z!�c�_�QEW��3(���W�:I�@�E�1Y='H�Fi3���ӛK�E��r�9z��4<�{��ڍV��5���!u������[!�Qyʵ��z�z�vPGi
,��S3#(��.~%|E?�ʆ�|Fj��ŨK�
q����ˮI
�4�RX]{Ԭ���>�#�;&,߹�Ǯ�$z��8ձn������C��#�c{�С��|��?Y��e�p݁�e�/����!�B2�w2^��C}sv�9f��@W����
��|��n�_���B�a~k�ƨU_.�W�TB1��w{��V���}ЈX��KH��I<<�t6t/-��xS�3' ��*X/|��D���t��Job�-�w�᎕l9���ۆ{��3�w쨭��?K���;�Ev%!_�=��B��ă��J��W�:FJ	S�Gypx��#�������O~���"%s�-Mn�y�y_�M����e��	�"$��5VB�<5�����T�^�uK�� ���j-���-3����۵�r�Q��b�1�mA���o6��'�y�(�DE�U8z�*2<�fl�Ll��"_O6�B��ʹX��C�UZYG�U�M���:j�����8�����.��¶v��._c�R"�xg�u�鞴M�s��(Z�Ѭ˵����m����{�0��g������7�A+��XU�^\ka�sKeh��51x�qk����:#���i��Wb�pv:<G$=����(�/i�J��hv�)0[��Wg��W�k�|1D|��ܐ7@5�0��t���t�#��
�����Kjʰu�ߍ���;�W�]�b).�P%,�®����V��d��Z�σN�awK�TO:)�H��}g�ȈT9W����PTk d��+�g��9���9<�dSR��35���^ܼi����ް��Ũ�y�����4��,���?��]������] k��Rmֲ"�wt��EZJ@uϢ��`x�6k�F���9z^~-?/Ɇ�
���̡G�����zL�_u�����댣�Y���{�ĭ�B�>�Q��=Gk���l^�<U�P��k�`ޣ%����������vV�1�Zл�>D9��a���({�l
P�l�KW/�l� �6C���'e.\�ݐJ������|u�N��饾m��i��D?{;%A�;#��&:rYs���В���Oȶ����]%΋ ���'|��޲hh)��j�:k�c��f��<Z�)�!��8�8���m�r��u�%�o!�4�����%�j�����4ae.Ѷ��6[I�av�UpH��F2��F+^�%��j���Y���TI�_�*�)��������fR�C�e��HE����"�5���zԥ)��e����#���IW���ݦ%�M�W��IG�U	36��>���Q����y�NI[{G��:)�yt�|������*�A��=`��P܆g���r�]�b���DO�*:׸��b�2ec�=ZC-�8�3w_�̽R�G�ɫ�W�[`Π� r�ȅt�t��G��[���J�VK�O�uj�+m�cV�X^s��
`Oe�.�A���k/@Jed�8�!��ލ�T��J�D&�y[���]�r�����U��u�[9��l�M3p���yҶ�R,q��;�C�bi�����~�.^��Qf���P�׼������]�zJ�X���t5TX����c|0�6�ɏ��G�A��"A��^������V=� .��߫�B����2WY�
��l岎�CI�b��x��ݴ
�>1��-�������{���.j��?{:�}{�K��
g��=á��Jٚ�]��#n���e8�4y�rB����	��^�
�=V�%�2�
*(~����7��|���a~� ��=�W�Ͽ���/}���{����E"Ԕㅌ�Ӗ���8��lл0-�� '7�"ׄ
�Tȱ�v�p��U��2���Ƶ���`����q�2�eIR��4�D'���
 #��z�7�'Ә�oh���oܓ�Y+Y]�	���nƳ3R�s<����[_��D�f@*#��j���dnу���L@i:��x�Q�^97F���������(k��1P����K>�E�������jF���\��Wv�}׼lE�*ZT{�Ǩ1�)�W#Zm�z�<�� �|W�V���u���YJ�Sk���5$ś�W�?�,W�=��<�1�9n�x�*� �r/u��u����]q�j|��Oh�y5�2%��Ek�����Iv|�$��ک4���u���b�����@ȑ�Izs̧�ep���-31#��! �͏���R��V�uQH~�Qr��ַ�H��-�)��{K.��@��Z�R���㱂Ar�肱�M���������m��y����Q
�����y�Ϗ�w��/����K���Z�K�W$eTi[��.����~/�h4�֟w�V�>B Ѽ�x�V�SI�.jw:Ey�׌c@?nZ6Gg٪�e�0Z3.�N�W�ݐ=��kҋn�<=��x�
�ΘWQ���a{J7d?��к�w�=>�������'A�1K��$��=�n�V��u�Nj��ފ��8,=w�MenQ�ý�����HR]��WYm -23La\L��,��%��MH$��3�����O|lx�{�	B0�m�����P�ax�/�� !�t@l3F)ڵ�j�x;z��n�2$��x\�^�� ���߳"!���(�b�Wͻ�y�m+�}g�����US��\@���:���J�֋^�V��@	xv��2�*)�Ne�3�l>����
N!hl���7^YS~/ec�q�P0�èxg��MMiQ Q���Nn&҂����^�K�YuM�窀����[�)+���j�J�;k��o�.���+S��ז{r����=�l����VYiy�Ω�[ՔݸU�������Elb��66��B�IM1����E)��a���SbxM�fK���A[""S1^�Hw�a���7��0��(�Ҁ�h[�iL���#v���W��rx*'�@X\{תUMO�g�ZQ��X5�W��
JZ�ܴ��ٷnc�D�N@ش� 7M��ē��֔EmϘr}jb���)��=Z�g��ޫ���j���Kn�@����r�	����p�X���8�k�ڿˡ����ۯ{��G~��o���'��ϔU�� G7q�Ȳ�w�':����S��,����Pt��.��<��9�JW��ʼJ}v�Z��ݒ�����楤�(���m�\rX�>��CV���<q���(��u�Lϧ�6*1IHS�\�~�1YO�x�^�����7}��|Fp�ŋ�$U�	~9�+�Q���:&��B2U/x#a�l@@
)_� ��鱨#VKj�j��-�tFJ	8o���M��]���E������	�y�y��O~�Ӕ�m^}�ᩧ�f0��&0�rO��q��-���T膱+�Hge��7���q*T�9�x�h4���_R0�KB������s��R�׬�@�[�,�v9�z�Ƭ�o��wc�tLq�e�nb4�jVeC֓�!<v�7�w֫�+���c��ެ��I�t\n�n֓��+��<���n|�=�=��yo��e77i�+�3^S�����GԸ:FO
]B����W�\�cm/f���n��%#
��A����B��Q4|R V�s��)���U�P�0��
bI��j�M�����0Ÿ��@�9
�F?R[�����9*2_�������%Rs2�z�o�O�u2
<`���Z�;E�8�m�\��kF�
8+��ll�o�p����G�40*�P��Nm�y:kc�h��e�)�kQ���k��9�~t$A�Ǽ�fER�g./��������ܦf�u���n�%~�?�(��Ɠ���o��O~����εw�
�mM��O�K!���n���&\v����=,>������r���ѫyLSAjn�z7�S�h� y��D�aK0G�E���jy�,��N��j�7=��5�^w��%�J!�ICZ��$�p���s͎9}�\@*ָ��>O�tۢj�Oר��f<�^�8U��e�w�<��)�cJ����ޞ�VaƉ����Q��W�x��p��iBㄉ)?9:i8��+
�+��u0�{�9�Co��Y 
�e�����KW��g�l��:k�>Fu`���=�ha�H���$ż�B�:�fg�����&-��Y0b��3>�ɉ�]θ�<�z�`��I�2��LI$j�D0����;�@�}>��5g��)8}����S�8������K ���L�b�U� �8�\]Wr�^7�3*�������`��)k]�6��O�p�S�Ѱ��2�F#i�8v�b�����V�W�T��徎����;�jc��*��h�����^���ⶣ�y�l�^��,O��*%F�>3��ܯ�o�3ctdl�0�deT�'��r�P��!�=�$+C�s���|?i(17��ƍi���:p"L	K�U]m��Ϥ[7�X�ф�yp �)j[>n���^l�`�#�m���^�p���]7&�]�ʯ@K���*�3�\��9͚�TH����&�Z��I�*��xk���7���ٗe�u�wj�5O=w��#A� 	��Hɑ,ڎ�ر�(�Z�W����%oN^����!��Ȗ5��(J�8�	�����y�y���|>{�SU���$f�]`��{������w��8�~�?S�a��7Pָ�MGLL�v�'{�;8Ws���_8�.��.=v��O<��^�I�r�iC+Nc������gs��{UH]�In�X>��Ra�`���eБq�ߏ*���ռ���11�AxP��ī��JoR��5D�H���n��Nh	���	�<�!�:UH��t��aN5	AG�t?1N,��_uPlf����֙�����|t= ��M{��(��o}zz�����(t����x�ާ9�������`�" ���qOӄ�O��b��&d5r���	�,	oI�e�5��͓�C!7������dx�E�t��s�}9:�eD��
��e-]�2��z-r���t �a�<K�B=���~T&��ғ��zD�v�pI��=nz9b ���ǈ'�/#&�Z�'l�����
�\y��K!��3R���Cm�;�>��6I�Mf�x��Di�h��8K������ @�%!�#�.�>P�]N��^��=�w�2���	�vjl׹��$����iNg|w���~"SIATi���9�N����?YϞ�^�=�)o��3M����|�^ON���&n������om�9�y�J\E)��h�x9������{��l�׾�$�ͣI�/���
��Ԅ���=�1B��h�#fp�!�f<��D���(��c�mD<2�������*�#	{D����� EZ��=D'H�"*�L)h\YZ��Kܞcq�b�rL�mD����8ׂ	YȵiL����ަ5����w�R9�FI� hRcZʎN{ �ďr�I!�ւ���=w|��B*t�������w��ݿK�����z��<�N�hݛ�R�_g�wT�S]G�7�^���oGO�E:^���*��b��ӷ̹��[�Cc:A�G���BID�7`��M��m����� -�0P2^vH�SQ��^��K-��c�x^
B�#߾�n�GMٽ�����[�6[�k��ff�bn����m�0�ܻ)n}�fl�a�B����/ޖ�o~�s.��i��4߼�$�5<�ȹ������g�����m����7���w�ſi�,Fx�����[X^��:}�/##�51�NR�*���R&?�gM��5������_��*�4>�/��W1,|�Q��Q+N|m<��*<��Fl���]�G�ߵ8��C/x~&L�قYld�#�����̅�"Sچ�����4��^��|vP%�k4K��z�B���I�"��������w��tC�f��b�>�X�_�܈�5�=��)��}��#L����k�e��+a�1��s�~�s�]ĵEt ���;�	����{��Q�g�|6Q���y��O@�%,���\v����D���W|�Y\�on��sf��YE�A�摪�#��ܼw�=�1Ҵ%�-k#E�ͣ�H��d���M����!���:rī%`��`��p���O|�FK��
=B	���@�}@ӢlqluG�~z��s��*W�Ja�V �o��i�\�F,�tn���F�%r����ҍ���m�p����p��zpW�D�
��4k�p��l�\;���R����_�̧?��_|���k͘j
F�q+�:�"�ruq�� �E��S~?���Xy�.����R��Qk�;g'�қ,)��@P�����p����E�r��k9����w�d���8Ɣ�P�{X��O|2����nld%sv��h0i#	B� ?���;�34�ѪwF�!x�D�s�3��ͽU����ݏb��m!�ז�>=�wwP�F�<c4Pio#�`�����������e��fh�SF^�F��������y�=J�h�y���S�>�<���{��a�S6G=��[K�����f��x�/�I�Hң34m+�"������3:�Jo��P8P1:҆QYg��e|�Y�����mg;�"I���m�S�a0{kgiZ����2�c=�.�N}�R�ʳr̤�0E��������A3�ۆ�U��"�h��$�\��k�	��Ur��Y�$4������iC���Q{�3&�ah�y0,�*m�w��\�^z-�P�i�vFa�{��J���!�H[D�?�;���z?�9k�� ��<K��|�:c����6��:�9�Uʫ<��ʇ��MQ����Ƕ��Pj�?��盿���As���w~�f���!��|�f���g�ɕ���7����4	.D����U�q�{�E�u���>װ�g��OC����͘q*��j�l,�I�ݧG{C鵻�$�EU{~8�����q�<�����"�(�Ѿ�9.�=ƿ������T�t��r�������C����6�Cw�9ʚ0�GF���L�c����Q�������޹�Η)�z6-eQZ� �X(��ܝ�3��b�M�  :O�g����zj���G�~4��{�ߏ��'?6*�I��3o������Z/�56�^[��Q!9X#�z���� �������z�,r4j �������ߧ޲�<��#��_jVP��^~�ы���w�!Źs����6|�@��K|�M�'���b�k}����-��Q��?�'�L�4���Av������wx�4A*��ƕ���7�n�^�_��fk��/|�����o7�;�,o��L���~���?�v<[7�ʧ�e��yq�z*�܍��}��ƂҊjy��9�p���X��7��w)nOj\i�v�IU;�$���G�l�
+j�go���ni��K�>�]�a�D>X>�$�/\OˈI*9�~��n�$3�u�S��D5�H<�	�����>
ì�Y~��i׻ޤü�óm��#�z���o1��Wǌ�k�N���E�'1-�B�p�Qw$Y�%��}ֱY���f3݊W^G����|w�+hSU�W�!��f�6��ڴ�!�k	c��"#}���C9��V�ȝ�Q�L��n�|oǶ�e�V�s��G�n�.R-2��GJ*�0i܊Ib��8��탧�@�L��*cֹg�!¬�Ñx�c��b�H�tI�4ܝ��\1��p14㕩^��Zq�� �M�E:#y)��E7�s�^�����ǲ����]�/GbfDF*��d$G������B��|�"�N��k������7�L�\~�М�����<��u�5Q
�`�����j��͛W�����������,��\��W���*�����b�g_K�4�8��1:��z�H1.�nPDw�N�t�Bl��u�������M�ކ/����γ���S��Q"��Vtk�dC�ױ}Ӓ>,�jC�Zˎ���6�G}N����n)���ԙ�a+�G.>�<F}�Y���k�gt��SgC@=X�n��v��H֭��lDH/�1!�z�a��/\8�����͝[6��4�y��aA>>JN������w�S_v5���B��޿����1emO7���'�'��c�P�2B�
+��a�C�J�P0o#W� ����9�
�}��-��!L���x.
#�:�|�B3��:'~e�6Nw�0�{�s�#qy��x�o�8�����1#<1U��P���u����q��p^c�-���vJ�I�==,יU �B�㤰F>S~0jԡ����#��W$!��Tg�Do����фH�ۥϞ���7�RD��i<��u!`�U�������du[B7�z���;�u{;r��B�������E��Ѽy�=L�������q�vv˞���x���"?g�(�ߧ�g"��xQ�WK���g۬�m,��ք^���n�V]Z_l���+�{�7�i�Y���"�z����Vי�
rr�`�
�XnYFe4"$���yn$ͽ��*�`���q���xSWØ{�^	m	�4�����n��`��H%���(�רlG�O&"��Qޚ�6��=}Z���%Ⱥ�H/D�Q���#a$�����5<Ԝ\ȱ�+�c�H��I'�8����с^o���J�\�����ԩ[���g��G����>�~��]غ�LB@�J��=�\}��&鄥Ū,�)�±��b�U�'�CO��ֈ���?�u���+G��]K����#%�?#X(�<#�IC}w�kO�5�2�^KE豣�*����襴�?�GX�=��[���%�p>sU*�ȡ�8y�Ts�q�
�S�<�,�>ǆ�5F����杫7���o�e��ɨg6��W7ќ<s�cΠ�7�w߹�b_aR�B�����:�uȆG��$��������.9�7�4��/7����?�̟:ռ}��8���y֎��
;1�, �h\k�M��4� �О�����'k��4��)L��,+�^�k(t��my;J=��(��V�����l*�\j��x��3���ꈃ�u�����K/k���!	I-�:(��7���i����0�l�bL�G#��X��kǝ�P�~�5l2,�sJ#4�D&�(��ni
.K�_7l:��}�����l\��慳�B�b�HI�V�����_�ͱ��[�/�.�q7׼��G��`m�oɆC^��k�kP˥M�gɱ3�`�adb�Z&{�J�������o�ܻC_vHj�]��
ē7JC�gs�~c����z3C�e�����(�h�yWW�ھyg����f����� L(�rd�^��lf���}��"<����>�� =�>	��6%�q%C>d�F�'øK�Q�j�x���0�N�e������B�{�T����Jz��T���%�HDo�g��C�9N	��T��|�4��[4�Ʊ��Z������x�S���G�x
B9�G
�&G�y�Ԃ��w�1��/؟�	��ӵ�׺�kחZq�%z���ɯ���Ʌ�}����s���x~�ŭ7� �����*i��¢C�
E�Ǉ��\b~���BG�4B���������V�l�}XcnyH�F;�P!�h����rRkz�ȟ�?�k��g�u�_�淛7��l��2���̏����^�����Rs�)n��a��_~�����C(���:P���ϝk��o�6-gO7������?�I��dS{� ��{-<�1�(�Uo�� X�#4y�� B-V�THj2��>��%�>�T�)��d<�x̆+�#ސJc�TũS'�ڲ�W;����r���9C�wQO�^|�;C�[?�)�%_j�@�lݿ�A�x9��}u7"��]�B�1v�#��g�G�x�<G�s ���  v��s'¨[�q#�6�"�>��J4R	��P�vޱ���;6�!���-�3�����9�8�֜��~��Ј�[hD9b�m��kg�DH��Bm��S.]W�a~\�=�����`�5I�������ޛ?{����:d�:�ha� T:�z@Z�އ 	F!�LS��co8�O`��i�Djc7Z�F8-�/U`|.T#���s�w�hʴ��ua�Cb���о�=�H��k�p&�so�h�`��V�����b�raa��S��{�0z�ʹ��0N:^�21�g�fHB�xA)sM��]��ht��6�Q�^�������}�1�K�:�B��1(�u�J�a"�`���pB��.^y�����"�{��_�6�?��k�~�������]�l���>3��!�T��3�jC��wܒ�R<�B<��2����w��5<z+����l޽����vm.P��EڒI����G/<��>ͰZ�b�}v{c ��� �dhSoh��h����~��<8�Q��>�C�PzI��l�"'ڇ��&�8���8��Ge��<x@o������揿�fMB�^o`��)���j�Y�q/f�!�c��U������	šQ�-���O����5�2B�Cd&��d���5jӱ�	��mHv#��� w�ݯ�"7ji�ރ�D�f�;s���KHC)]�C��]O(T�Y�U�&�T��4���83�5(Reg����&N�a)U��a�!r\Sg��|W+�r�&q(�P��j�[$�E
�(�� �m�%�S>�K�K��YcLPo������f�u'�}vx>�[�N��ʅ}�-<�;����5
x�sv|�h\����B�����(0���@C KO��:�{Z���B��O�e�G�]���:��U���t$Q*J4S*?�Cq�U�;��hg�$��OC�&���Wa�߈5�VF�Qe���u��#�;�Ht��}Q���a�o�N��:��G�&Fnlȣ1���my���*� ^{�`��j�^��9�{G%�1u���s�F�H�3�uGe��&�7׉�i � 7��	+����^:�O�� ��'�ӈA8)V"P���:���S��P�g)������qF�P1z8�B��gѓ�)�B:#X���q��,t��/���	�_��^�r�%��]���2��x�D.=@Wwn�g�nT��RmI'0:X0��U�#.�x-?ߪ����ɼ���uJ�!uX���IH䷺\q�)z�FO��5_����^�\�jdW+-��|���l��?j�ܹ�ܼAv����L���<����m`1����M��k��\�4dv�]r�!��O�FA��n�o����|������uE%��A4 sz����;�|x�\�n3G�vgt���;ͭ{�x�vY�>ˣ�޻�^m���ퟆ���(�K�����;��_��P���9�����g���g����}ʯ�7�^G��	G�����2[+�՛��k/2���^�b�(�g���@�4�O���)��}��(� ��屍 d�?O�^G�)rMź���tJ,�8nx��HA��L��F2U�"	U>���m�=�����u����l�t@�7�t�{�����G�g?�k��T���aj�gK���	q��:���ll�JD+r��_�(���d7���gG�Ď�����dx��|��c�I~��6��� ���f�y��m�7�0IY|>���L��U�*i���H;6}'[܃]��h���p�I9aX����2*��D/u�ϝ�5�o���9���1��������s	4�~���W�������Ҡ�%63��|Ny�F*L1J2�y�vfA�T�4�k��2)�2��4]w��Ix2�E0��
V���K��*���&�D��{��{<�0���uי���b���N��i[5L�f�>�T�L`0j ������¹��'�z�&R�1�2�p�=;�L_��c%ω�C���Ɍ�#���,��m���˱P�M=x��7��k��������y
@i4ei�󈨻�)�?�uif�]*��Rb�l����pQx@��b�J+[+��t�o:噬���$�a�'f��^&(����{��6?iX]�#kWCXi���l ����L`�z*_ϣr��娤�̑�ם����A��y����8�ę(g��
Jr��,k�C�������^�.������懯�I�o�}� s�J��L��g�p͌��XgN7���f�HǹՕ��������!B��v��=[kd��\�cey�y��+�_���n�CڻuoeI�����C��B|�f��1��1�>��Q�-�7��<�(����͋W����9r�Y~�W���s�$��m*+{�'	�7e�ut�J�,�:H�2�e�s-�S��NC�F$z?]4I��)T�ڏ�e����1:֫1��"τG�jTH�:s��fm����KЮ��LH��e���V�?���^��#z�����5w�>��k���������0i��w~��f��^ZZ�}e�ڻ�ܠaJ��w���j�S?��#AB��ԑ%f�*M�s�qϸ�:R��]��5��g��?{��5����f���WY���	l~�8��'��x�\L{��p�z�5B�o�%N��_�00�������D�a���p�^�לY1�֘JْJ;����gg�rQ�΄)�|p���������Kqh�z_��4�n��e�ӧ�6��?����=������i8�ϟ�K���v�OK���x�x�^Í�Q�K\[�jr��I�����M��ɺ_�T��{8)D
&g��i�T3C���g�O�;s�Tsc�k�����	h�2��n��2��([;v_�B��T._���/��7>����<xx6C�.��=�p�1�<��Oi�f�N.�͎�SX��:e�לy��m�;B�~�ͭu��2��q��F�cR��P��zZ�Z�6����^�~�T�%S\�z:vO2g�ʜ��dBieu-z�v��h�pax
US)��?w�酱�5��y��K<ћҫX��jum��x�=���Rs�@(����F��!��qz��d��$��� [83�d3M�{����I�+�<N�׏��>z3ؿ�Ԑڅ.zr���̟C��Pbޥǟhnߺ�ܿw�&�o��+��Լ��_n����Z�n���%/��ֱ���E�Y�te|�ĮP��1��i=̃��2�>�f댍�I]�#�RqxHԷ/���A@����ٍR�w�y��6Q��a���(]#��w�}�XV�|�\����d�HG*�n�)���i	��>3��9P��	p(����jDo��9��<�B��
��e�U��Jɘl�0�r����r���Ϝ{Kv4�3��<q�D*#PAZ��W�i	��R�<�%�,E�{�V���~q��ѣnB��;���;�M�"okԣ�/ǈ0|��7ud����Wx�m�,��R)g(7Yb��ez�ɺv���+��c�l��KD�%ԙ>ED&�[C�w��r:��yD:�VUY!G8a�a��Q�x���ᣑ:��VXx��v�k<Rg�y�1.���d���>�>���+ݐ�U"\�H��&Mj\�aH�~���z���ݨ�Q�q�;��p��L�<��M̳/�U ����BD�B�[��
��������K#�M� �/s��9"Xܛ2��F�~�Ȯ�P.R\���S����C�7����� ��[�Bu=��\�����<���Sa�u��a�4mشP;�̕���m^8_3\G�Q0F��uu:F�cG�;�}j 
l�˭G����~�f�����)�]�6���V��I��b�Jx�9ElOp�\�3O?��C����u��z����*ђ��@�4'��W�D-�<�;`P�*����+���[�����?|=�h��]{�5S!$�Cs=lę�y�n'���#�t��50�18��ﾌR��&]������`���A����Y�;��
V��o��5�׿�����|���@����y���w߿׼sa2D�{��5����(�9���fԟlk6�<+�(r�>���!O���G��4�j���k1��0r|j���Ț^hz�9���O�A���b����8^�]��٪�<���p�^�2]�T
��7z�%"��hg4 	R�%� 	-��Q��Z�t�g�Q0���}�{��#ͅ˟h�=�l���?͜���'Ϲ�46�5Ԇ�e�o�[�pm���� �E�kX�~��ݸ�u��p7�\Lb�84���C^3Jś_Y������@�ͧ�����z ��2Jѱ�;%Fl4pɰ��%���a`���G�Bt-����:�Z���.�֥	BF$cr]>փ�����fWF�,i�Gh\��>��@�U�ǕJ*�x�i�E�O���;ʓ�Bf�|��}�s}v�z��4Gߦ��|�aı��дL��9����tc�� 7�v�<,�nu��<FZGtd,������h`-p�K��V	��qQ�%)�S]���e��F��0����ĵ�^��V�3$�R:E��)I�C��SA<��d���~C6�>L�}�e�ܧ|l<to��ŋ��~��~��_�Z<�8�lx6�;��Ps�-��"��B$�L��.��,H���>��[!����IO�:!�5$r�V
.[wZ�)�� ��W~�|�s��1=^3Y�d����M�Q�x����{X����_~�2F����;������fS�v�^�ܴ��fJˉT*���*pC��~��#��ؼ�d�oSC��z�ܬN\�%to���ר5�<nn�c�Ż��^Bl4'榸�G��r���*�lj� K�����=��3͕w�mΝ=�s�^����{�o��5�8H�e.?J�ރ�F�ʞC��%����+b����WX�5����_d^�B�7y�C	�$��ģO0��"���Tx�
l�y���De���yd���l�3����g���n���L�c
�%BZ��7u�A%q�4Ó�2��������mv���-y*�+:�+:�2\�M��z�������Dֿ��Ƹ&0P�R�{�TP�<����xt�
�4@�gT!��S�������R��׽�Cś*��a�λ�4���ꗰ|p��s�M�!��?e��+ �x,���WǛ	���Vct�t�h�t��e����}�?Ԗ���i~���"��r.2]l�ċ�l�2�3ܧ�Cy�z(�}�ʠ�@n#��������2U�Ai@���5B	e����G7�Svz�"i9;E��v`�X>i�M#F��&?}�1�V��ȁ��.\� �'$@��oY�*�SPF-��*�`�aǽ<|�u�����PNd����Y��싈���x�� ۩nxx࿟�{��t�:�m��q�'����WSo��7=�����d\�*�С��J6��V���v�ux	*��g��usG����J�dj����z1Q��.�6�/�oWu�BE���[��zv8�#BV��	)�}S(�	6�ֿ�H�q� a��^��g�m~�!�0�/.�n�U��LY"�72���dS�QdG0-e�7���3��M���V��«�ԃKg�s�ᙛ�X���U(]-x=G����Z��f��Vs���4׮��\��Ǧ"�֯�V<Ke6׷��$��=�pq%�1�}�3��O?Ƈe-'����[5���]�C����pvi�s5�N|,�'�m��6L9�2�����N�����X<i��?	>=��L���qbclj�9wz~��X��g=V���;B�5�^�8u��J�{�;����''�)��D=p�lF�3֖�\r��M8��7n���й旞{��9��߰r�.`D3Z/�[k��[���u�K�X���K��εJ4��?�l?�.%�Z72�Fv{�v������a^����&�f�8��!�{��y�q��zޡ{!�vI����;e�ʾ��7�Pm�U^~�[7��=sv[Ø�F<1�s�˸\�q��MິL�j�K��(Jk ��1�$�QV9e��DK0z���{�ܠ���<I7�F�v��Up:��c��9��JA�t��_{���0m��tEK��g�g�<��3���&����SZ�a�M�0"�٣unF`���1~�������Cw޹F����}Hwɓ�bX���  �I�1 v�$�=�G�!J}-��8ǡ5�>����X)tD��/����޹����=>;�q,�֒K?pi�����R�.sS�rm=����Q���!�k919���:F�	��Ó�i��9rz�i)j��nQ! �[
��)7!���G7��v��<TԽ���;F/�GR�,�M�a?�$��J���tu{��w����:����}ɦ"��� ��\���"tsS�}��5��&�-1eM�������r�+^�fQF���ԓ�4/>����1�2���W_��N^>�O�[O��l�;�V����|��Q�x��K�����ʗ_ʦ74�09��z���W�`hc�)]>2��6B/�A��yB pQ��B��SA�:D?�2�%� ���)��I����`=L�6�?~�R��(��òw`�^^�
��O�z��G��g�'5���x7mM���T�l�ȋ��_��F�����x��k�B������O=E��ts��"��&7	%�`RC{�-��]��0V��(u�9���1��v��*�Nٶ��S�b۫��?��[�|8�ۧ���(��?gX��y�qE*��g�7��"�B�]��gv��$��?4<~��ɳ��bDmӼrx*��T��5��=n��T2�Y�7pa�u`~~��Xo*F+7\�A���ޛ�$���`�1�'�6kr)B~�b�=)���12�b������H�$J��1>9D��0������$G���z\���i�|�:\�&[=�,䤄R۷���u�~�a�G(��u#��ǝ����`��q㔌ҋ�	k6��=��Ĝc�u�:^��իW��~���X�_�9�y܆)%Z��	fy*��n[/$���e쯻��⏥�v��nY!"�Y�VTt:>Cr*�l�ϼp�k���gb�e�z�a�g�~��C�|��]�ܧK�|,�Y�鲟͓����UX����-���S |�l��~ȆԚ=�dB��6�2��R׋��V(�$
z͹�N��{W k��;W��5���G����wjDq-*!�q�(|�<���&����Õfx�Q�\�]��3ǟ���bJ�|yy����#?��o�Ҽ~��T�j��_iN/�i�]��b��UrJ�lQú�@5W�Ad6ro<?���l���<d�g�>�H\3
�V@)��w:%r�H�P�fs��у�p�')���eY]�յ�ם^ZF�|�3fb"�zy=��������R������!��^����w����/�����K`u�����J_>��
��O]���//�u��ur��r��YD�O��`���&�>��,�>�A��x�u�@(i��ID=���Ͽyd�S��;�����ȏ>���M(Ep���"�5w���5��!.�h��k�����ll�ޱ��s�-��Jn��GK���ƥX�pA�8at�e�.�=r�`;Ȅ���r9�{��T��d(���!�q�^v�-��<q�L3-�ޒ� ����!Ah;��C�є��K��e�|�K�n���u���r��ȑ�,/Dއ�U��<�I���{"���0�|��gX�}~_#�O�܍��"�v��^%�؃O�\��#5�5;���8�7u���W��/�����g6��';�\&q�&n���G!OR��`�=�r�a�Oi�ƶK���T��26Y����w��<�DZ�q���fX��
�ŮG�z&q]�����s�����i�q�����瞍\���uk��{�)N��ajx��o[�v���t	��>����GH7�Ru�VO6s���P ĿTT�d%�HV��`����L�a�u�@�����/��4�hhX�Iәw�C��z��m����(���?l6Q��u�p��vg��à%g��t�ù�����fh�^�D��;w���u�I28�Լ��¹-��")�1lM�����|L�B��Y2h�,C�v����;����ľ�A$rB�`>!N��<������4�7�8Ƣ���ǰ�9n�F���$I�kc�)��Mmvv��=u�9�~�d�"�L�����2Z��>C�^*B�>��\ �#���|�`D�Z'��_a��T�"�z���kD:iU:3����OC B�]��#��`�yu��܅�;�h�������M~��G�]���l��������z�t�uQ8��ѿu��)�X&�%��իH��,��n� �����|(Cd�GJ�Tp �_tW�?��w�fɛQ�7����������$��p�����8��zO ���'��GY�VHl�������4���}+64��c"���Q(�_͡��]p	>͚S�dv A9?�|{�K@�;5r*�Y�����G�6鸧w�	���.5��§��g.`���,S\c���&��0�#�M�1ׁ�J��1#'m���?�������[o���7���������G_�vwz�~��vdX�Ji7R�M�OJ���(�|w*��ׅ���R�'9UEg������nkSUzZ��o���N��>m�Q7��,����G?mN�3�܋�b����h��v��Azb�tĩ ����c7�?A�°w��1Bɩ��v�2���|t���q���k�L�<u:Y�[���#�^��<��q�Q=K7�����|^k���^�*��k[�ܳ!���y6�F�����벱���G8|}e�z7l�E~��[;\����c��$�-�J^�Q�`G���x�He�]�8�)��#�w����\���JE�W7����!�%�s��Ǔ��j�4���d��g������o�x���O~�q�@�EHv��=��pNC�>'��(,���n��m����\�Ao���7���g�ˏ_�S���o."�ei���9~r�m�!�G~��m�v|�*�a�ƙۻL����M0M���Ge]�r�Ր�Ǿn�����so�������+���h�'��{0�v��%F�/��G�w��Q������G޽�{=<�xV��������N4��$�m�0�YEA��0�c�˨Lx��%.<y�Z���4J1A�������tOtf�c�8~o�tK]�T�7Fk�W��M�������.uhl���`s��4jb*�r�ՙ�8OCsxġ497b��Z1�4�nkVz7�u�c��vpxtbj�ejl�-�d��ټN���g�w6����4����^��j������0��b�l��Ϭ�_�_����Cy����k��O�x�3����c�A��r�k(�옵C�h�j:7Y(:7d�@���h��ôb�l�����6�B��:1&�K��[�Ӑ��KS���(��gRK]'{]�<��6�֛��A7�w�4�.]���s�Vay��nR?��՛��Ս����ۥZ  HUIDAT�]KچCs E��ƹm$C���6�a�g��i�)���'QGJ�v���åuڪ���;����v�G�a�b0�������^]�)�3j�ǨR%X2���[G:Ӝ=�u�����8�@#�.u}��J�c8�k�)o�(s�Y�gas�*	���n
�s���G��e�*N�N�Q����K�)�i*��	@��eʆ�	�0~����`��S��������,�O��g���\|�R�s�!sb�1^a����
&��5�W\��g8��zΊ�x=S��kع�F�N�7kͳ7=��f�Ju�F2��=h���5�L�"���Ŭ�e�w�4s��{܊���`��rnR�/j�s�v2��*ǣB3��ҋ�m(,l*��R���7�$�U�g���{}��������	G�L�w{��Н�{��U����z�aZFz'Y�9�������vWf*/'��?FYbx�F�|W�F�"�qzvz�Ү{��d����F��N�M��E�����he�;91��n�H�͕OQ�Q��k� ����=��<�ϣg���5�ǭ��'k̓+D�Q���������%/��t�SO?�l�
��I���^�~��$�v�}�`r���w��${f��2gf���~����B�+��o���W~�W��������(�q��a\E
D?&��G������q#�s��ݒubr��0d�anM��XLU�Z_��[OU��e%t
9��ءl���"��µ�a�|���Wv����{��w�����c4�җ�D���[��х.�Ʈ;��H��IbO�X�2Iݘ�a8�G�R��Y���2�C�/>�x��~�y���j��g��^�&�,�y���u���lR'J� %�XC��1��k�������v�2�l��2�9��BIwc�Y��w��H�FmXh���c�q6a��:vi�3���/��1I���Q���|tTNvW�Y:ųرL(�xX�U>�K�)Y��+N��v��`R�����8?�vn�k�k�u�`��>����Qϫ�Z���{���U�P�a9�Ŧ�Vb�_Fc�ퟎ1��������Jz�b��t��:�W��lךs�(7%2��8,a����T�rLI���ڟ5�}S6��s����-¤��#Y�1"n�1b	v��4��mj���q|��c����o�1�����|6y��{Z�m�����������ͣ�L�V�`aF����n�%�BN��B�9��� ��8=���ud��q6�r��>.q��=��x�s��S��)��ӡ{��2��J�,Isg���)����V~��"�#;�g�-y:���%7'K	^7��mSNe�ۻ���Pf��ȥ+��,-^M��5�,=�ه��P����q��%���dD�8n�N�7o�n>�y����2�떽i�sO\���n��I��5�FPE	ɱ�:�
�'u�ɧ�����o�ӥ����/���כ����6t!��UٹI�D���Ʌ��f��Hc��ް��4&!p�N���.��b��<q��Y���e��d����܃R.�PZ�jT���%C�2�������9m����4�Ce�h?�*����ߣ����L���"��%l�0J��B ���G�"7o�Bq,E�n{�u��)��d��4��ܿ���� �G�J2��KO�Y>�\�v�9�7��M�g�w��3of_k矽�w���X!Ң��� ��p��L#xْf��ϜXEvor���k�lO쟊����)>$����>�`�}l����¢]G���Q�J_3�s ���!?ϧ(1Ϟchu�ڔ���Tv�`�~�l�=�V#�����U� c�ǀ�qs������~2	�zi��-+��w��j��=*$"�ӯ�����Mw ���K�A\D8��C�� �~��t��ˡ��k�\�:]��Xt#���ꆸ���t#�_��:ls;F1) x�ܷ}�!�]�+>�9�_�|8:�U��NH5�s��r�=����:��l�%�ށsX(y�~.���EW%�$hp�H㮍C��{pww����� �!H���ڸ$�;�7�������թ�=���s�V�����Y����E]׎�@b�׊�]���xog5J���ߔ.��!��x��������<=�&�Ȕ���˅�u�MҘt�I���Į��_���n���n�\��)~�p�~:��2o_��w��s�<��"a�iv<E��kO*:^NoE�w��⾸g�F�`ҭ�
����U�a;I9aճ�G Kl�}M�S�5��ou�g�= �I4b�e�Mv��%���#�<�ȭ�
Q㺞}hQ�ԩT�0��f�Zn�x=��5�T��� v}ZǍ=~a'�<;�F �ɂ��7���� �*�`���Roj�NJW�Iz�W�x+�V:t�S��Nlj����⪝ ͚�m���ڙ��B�hL�.�儊PK܋���G�9{v~4�&{�3�ݸ4�:W��*�+�o��8ӋR����q6{�L��J���)Ͷ1B6��!���I��e[u�g�v�p	�J0�`��0E�JF�B梠��n�O�ȷ�o��"q����*�H����m�/*]֔����8$�u�j�=-��Ƈ��w��`���ˏ��q]b��I}yΩK�pJ[���<�/�$��_��E$;�aKN�-aKN��&��Drrrh�=�P���Nĺ�U$O�G+��Poq(PCŭ����Ϥ\6)#>n�K�0��1b%e/BW��U�4B�#��k"��e���+�.^�E���T����ާة?�6MZ�������㢶�I��3�m��'�;=N_���8?+����%���t�jcK���A�-��
IDC�]K��(7b�?�����~-��M�r8Hز�E�?�^O�ǹ�H��:w���y��S�Kн�5w_��W��H<E�g�=�x|����S����t�v[��şQ*/_K��D��(�~~�u0�����u�
�LFȰ"i��l��p����k�p��<�Eq"��;4�
nI�=,�(�qm��|$�L��!㽒� ��E���=��~t 9C*F�{�nOcCs%��L��\��|��h��2�(��J��g�J��mE��ց��h@g��;b�Jy <����-W���6�y5��A_殾�/�'-/n��������/��?-�a>,��H��X�����Z�5�	��c�w�fhkw�R_O��2�6�$���mʲ)�]�>���6�����]'���\����/�D=����Q�LD�&�����8��mG9މ{ަ�/��B~���|�f�
���uSc��w�k�@�q�N���&����e����Э��(�����71C<�� ������o����Asu����s�ߐ�-C�[�c�LG3R޶(��y�����H�~C=E|�}.q�w'v���6�n�-5a�QS�m�����������ƀ�K�GLB�<�˔��"�zף���w�����E��w��c�D/�Aa
����~9��6��?9K�G&�$�H��2I,��4��ծ%�c��{�R"�g�� �5�lfy�V)��59�Y9�w��A��1��1s���Y4Bu����F�\�-��FBt@��bz�֦�p����aZqy� �?�\�R�ꯌvwٶr*Lv�s��Ǌ(�ħ�4=W�8�j���K�$B�flٖ)t����0�*���L!5��W�w.� �i���V�X΀�{�\&%!�},�K�}���MX�B�駅R������>��.��K�Uw/�x���f������7�d���ͤ���l���ø�p��:ŔX��@���/�d��������;<�i�}���:m,��~a�.�H�����ox�������woA�����<�1ғ��Vγ=���>�L\�x!^�Ͷ�<�4�e-�2(│�����?v�a;+����Xt����Jç	]�H�l�&��q�͛����@Z����[;X��KS���������Y��@�D�'���!v�M������#7H�������<��\�����{�J|�������6L͡�������-���E�KjC�g�A��V0E�oc�ݍS��>�Dx��{� =*l���kd1���A����D�>�u�+>�͗�ud?��=�[$��d`�4�U��Cy|�%���$?��Rr�8uXDޣ����k�"O�a�"��`d{|UX��4�����T)��vCO��{�Qf�Z\t�WJ���q�*I|�򟍸h	���_�~�����%\����})�Ϟ(�bqsB^���	����J��s�R����M3����ޕ�׋r�����V�L��zʄ��Ϧ�ĸ_��"a��<��o@�v��ߵgu;�L2k�c��n^>�(����S���N�"�}6�?�������f�ݚ�?��H�PSf՗�k���Z�W_(���W���>�i$�M/dA=�����	;���O784�H0��t���8�"q���#�Z�ʐ�1�F�E�^�R��)�����:�Nh1����ۚ��}&�֚
��0��ڋ��R\E��ܞ�h��y;/yZ��X�N��L蜤=����.�8�FJe��d~�}��&H����7ZGϏ��/��uX������v�&f���Qwn)�^0��w������	5�5�4ٱ������vV����^M��1rظ!gQ2ć�A��h�d��'��d��r@��W�����V7�i��c�(�,������橷��j�x�<�a��_t�E	���>�&�82���ܚ��R.+̳��8Vɾ��?IH�^_X���Ą��]��;��V�%4�4'��٥�S����d���
��I	Y���(2t�� �Y���A:sp8[��?N�zs2��/�E?l�Q��srS���?@JϢH���S���pC�U�36�e�����I��%��+j�XJ>�)C�5!Y����}SQ��nA��s��T��L=��`�3����1^��A��)���-}��"Y
����b����Z�nz�+k�DB:#v	ݓ����r)��P�����0��.Hc�Yu���S>4�W��5�$$�;i�J�Y���ß�&1'��B�Z6M��T��?Q�Z	��yE��0Mk��4l��=�V�ߎZ�з�cu�-�3�HbC3����ihB���d&���	�(��w�g����,�?�O> �v�E1(�#q������R��J�?!-X�Ǻ�o �l7߶U��=�H��]�ϛީ���2yP3@p����:z���Yч"�@̬Pz����|I9P��bvFԢL���c�H]�)M�Uq���_��y`��.�i�#]^X�[�*��V��eh�BEn��[!���SY5~�j\	�v���.l�,Mk��>_F�ګ��8�<���8� R<e���bC5@�t��ň����|xa�CdS'��-��5���q�Z�x�=��u�w�#F#�w�fp��ߢ0��i�z���f��]Z~�s{p�e��pou����F"8��CT[�5�����'=��WJ�9�*��h�l�~��BD��G/����-ŝ��D��=jX_iD)��;SW�bt%��2�l�.�_�"S���c4�uJ������إ��v�Ć2�lW���1.L>L�:�l̪P�%����@�/�US/A�1�%0D���	Ks�^����AI/#��U.r��v�=�N�����>�Q	��k��4L��-�w9q���9QfŇcg[no�Έ������U&�rm�lə���9y ؇j4��(�oY���Q�y��kŌp�+���B{�����C��q �� .�K�"����6*I�Z����[�ka�W�^��W��7E_��r����?�m���|y���8�>����no��O�%?#�l�u����6!?�k���!��[�e���438��Y(+]Q�9ñ~C=�௜�#.��p�o�/Y`�3��4z����,�o��nBT���4֙���?��B�Oa	�2T�pL���Q�F��~x���凜�+���&�'@��-�I�D®I�B�I�D���Iq���X��@zy6�G�W2L�~x�V$8'�v�?�쐪XB�#|��︧��KB�OI5�0(96P�ϼ0�c�3{��rj��<Ve���!S�RW���;|�&{�, ������@Sr�)��[(2o��&��w��_BdzH���k�j*2^	
n����?�A���	�������7{_�O(����k��J�@]g�����I|�� 4�u6����'�D��G~u�.�L`���3=�>>����r[pH���5�&�X3�ծ�=��A=p?yza����g��ח\��b�kw�}"ל�<ɞ��aMK���o0N��ϣ�.M��������#�.D�i��r��	���{�\�������゘ݯlx&��	���D����Ͳ�s3��T���EF��	W<�e���#5����c��[|��+߹[���#%Rm'y� ��I�ci�s����b|ܽո�5N1�*v��i��p4�������ƌp`�wyʹ+��ʒ���'4��۩���m*�+S�C�$��b�B�k�}��3Ơ���S��ϙ����N\)Jq���.�^�`$��Lwx^�_tŪ,����TJ�&˖�G��G��C������v����#����դ�-��kQ�ךy�A�$��N���N>�\���gwQ�&��k�8@W+�ػl�'�X��	��Kb;^oL��͹8eo�ocg:��c�ϑI��
d>�8hRDH;���$��{�o��9�<��Ta��p�)����������1�k�k��U�	!0�H�3 �3L�&��#�F�3o|���'���W����,.0bK���ҡ�OO\}#��F޷���,҇���F�Q���j����9�����eM���=�{;w�+b�;F�ht��&��
D�<�'N�e��j^Vk��ؿ�lw���q[*���.L8�[��]/t�-}��Sl`C�U�Sz̡7���<�;��O>nJmc��	���
ϳ	�&�T��2f�JH^=��w��:bj��V�����[ɌC�����Lk ��~�.1.�r�h�G#�Cg�	12|/�@�� )ة�]U��'s���>���y%V0mrm`އ��	�	��M7�6��u ��R�r������}�⯍�1�<�	 b�f��Ŕ�����P�Q�-vr��iذ
�d5�nɏvb��^2���Q���''Zہ;-���OO7t����@=�q��t(W�;�j�����	�� a�phDHEjl��"��_�G���;�!�ҊnzAh���@
�<iH"����Mn���s綌�B�?�R�э�$��=)�r�/�㙮��;¸x�e�[]c�D"��4����Pթ�}J�'�qYN,���$fߣJмD$�r�%JӶi���zH%�ē�$�e�к(JW�ݩ��(?�Z[�P��R���y�$�f��3��a[�?��_ŵ�)[����ET�����_���\�C���
H_Ie��ֿa�Ji�����D6��I�mQ�m���rgM�=�)���	/6?ӄS8$ES��U�V�D�Ub���V&n�p1.�wxaP�+��,s�$��o^k��hBf/��"����M���!�5��O�l��	�j-���C�bҾȪ�s#���S�~��j��I��_8��uXPζpDYG��!�RFvKO���B�S��P�)�=Ձ��(Jиm'���iC9z��W�!V�vR^h91�zC�A��Vvj�V��/�7�!5������?��Y`Ʊ�3�\@�u霠(n��	�%�05?mǒm�w���|HF凭��i�m��Hu����2���{m�i!m�R����Ũ/ %a/@�G����A�T@��c����/��:��5ޗ��v�5���䝯�\^k��CWG\-�u6����7Q:B$E�x��,s�6��Gו�J�9zwX$$�A�ɥ��>��W]p��)��Q�)i%Qض��GG@paA��u�q�P�'��%`�9ٯTń���%�P��!�ݠ�(�~h7�
��SY8�,��}.��Y�e\-��{���M!8yb.��uƈ�p�z=@�Y��f,�R�&d@�A�E������v ~������)�u��+t���R��.9���+�$�M|j���-���`��a������k%t��;��Z*�8��5B)|Uh��ӕ�xM��?�(��aM$u6�����*�C��6�'�V�E�a�<�`�R�E�X�D���?!����R�[��b㎤ܔ�I��]3<�y������8�(�����大��c߂��il'M>��S�����5H�t�%��Cg���P��#����e.�\mJƏe��]&�gF�$4��Q���O�(�`����*h5ص �gt�Yr��X��XvnEk�rz�yW�\�P�/�G^��#���1�Y����N��;�OG2hUǬ��i�Ձ+��E�۟��]�`�R}��9�sgL�//�>.'��*ċG�1S�T�<5���F-�C^'��oF֧u�1ǥ��"L,���u�|H5sNI��� ]���P�<8=��<��ŗV�,3>���~�_
���{�!�g�)�ݬ�БIRLI��U�pĆ���@�鵯���Za��X'NǥUJ����O�]�r��Ai�2>��s�WJ*O��=v��0�oF����\�F!~�E�-�5I��*��ֿ�nK;vn�{�G�����[����*c�̢��|�ΰ�)R�[9 ��)z��|�k�a�Uy��.g{�;l�`>�T��vM����4z߿�g�/���7&%���r�_��U����M��c_p�E�Ǵ�I&���G�Im�WmϹ�b*&�	�P��Wʤ�'8u��
2@K?���]׃Uޢ�2+��q���2�k�!=a,��F���ut��OIvH>(����}�Nd���~&���I�Ęs�e��4�u��m�Y
mZ�}(n���)ީ�	�A���0ԯ�H0ZNUj��P[�V��ǣmd�:&ݡgC@�l��(�?�UT��[/���2GH��3/6���&�����;O�p��
�y���/2�싚CZ3s�u�M�?�d%�t�8��O��Mw�m�%��t|�,R?��FIA�8��_9�����dJ���a�v[#x��Ώ�u�*���U�9���I	x!	�f�ʩ�z�h�'��.���Hwr��� iD�<=����?��J9�i�����t]U��S�� UK�K��T件R8TE2O~�'�3
r��I���>$�V'��^;1!C�EY�Ƶj��c�ڽo��%��S�RhF�*e��t�Ŋ�����A�W��`�A���!���5���:+��h�~�!����ۛ~�Q���� �c)�`���3Č�S���_Ҍ�
���µҖE��e3(����^�6A��s��7�-�~z�B�W8^MLѻ�R*5y�07'#���s�*�9d��Aa���E�����U�xs��&�3�`�WE�����B<����]� �=��SE*.��K%��?��0GV���XmS�♪��%���
w瞉�AT������� �<�V�}VN��bDm��l�F۬8�����S5֛��7��T*qC����+��n�5
_X�^��f�&"=ҩ!P���gG����jl����M��c��a^�j���}s�sf-���l��̽��w� I�7rM���^m�/���x��#!�t���:�ˌ�Zǚw�xy�7��K�UnI����~��� 0�0�|/N��\e�vE�θ�-�:�)L�K���z4�=�5J�d��n�FxN��T�x!E��H��7ܟk��	���K�߰G�d�D
�;҇���⟥�aV�!��>�PJ@�����]=_Fy�vC�eD�.�5�,��DKq��GG�m��aQ�MR;#bfY��s"̳��=�b||�<�{'A�g�;*Kr+;ZR&>9lZ�
�Z�b�%:d�-=������c`"�,�{@9�:���1{��_�{P\{D2��2����ۂh+6PvI
�$YB�8��:��T�/�p�/�l2��A#��������.���-��c��^�E�}{���m]'k45�!fS2�О(���9���t��M�	&�ӊ� X:��%��<w�Z��*�JYJIL��rg ���Coŋ鲔��o
f����Dkld���Ҫyo�~JW��1[Y�[x?MêOl�oG���T�%��f�JUTP;��L >`�~����&R:�X ��~p����ǕeT&B��g�ѯ�ҫ	Ĳ�B��bB�b�xlNE9��pEͽ���eW��B�$�a\&X��휂��t~�^��uGBأ���'�M����_·�;���D�G�g�\i�\,��,h���*�1۵\LqW�ٷbn�z��3ԋ1�t�o��Jg�Pn���pŀ�A_J��1�.�q�}�$z�]k����ɧ�Z��!�`�$�1&͚�O�Q@���ƫ��I�+7��cvߤ�g��S�
�/�ye=�$��7wa�$!�UU)�?��[��j�_z��b=��\2�<�����MϺ�ӥM,�dO�x���x~�ʞa�N���=���L�ƝY��TU�#>Z��ä�\���;l����3������_�U������uZ���Zy@��w˅ǿ=�M+!\��O}FV?���[��k<����Ja:�p�����0�� ~Wt�{v#������l��&X���,�x�<�7��B89�Dm_�Y�$���k��'Ĳ��<�'6H������Ǡ���{��z;s�´�ρ~*΄]���O�isc��?�׺��A��A���	�e���ۓ-Ҷ�}}�Ž_��=��j(�AK-ܹO��?�=Yٿj!'��n7�>'E��6�e�!B%�V�B>[�:���������J���20cX+�>���hpXE��k('��!f���a6�m?��U�U�M�ww��W����C�G@�k�Rhɘ��T��-�ac-`e�-f$���-�4��)���FM�/V�!�g��"M���1��K���6f��L��ƾ���BWڛuA0��5��mqjy�;у�>��7�������TWryգؗ�|oA'�d�9�["ԟڱ�sс���)���1�B:�%D0	�㠈���� �tL�̒n�P>7'@O�<s|����чo��~t0P���-`
#�'ۭ乲)8?��^�<����������_�y��o.3u7=%��7��أ:`��X������L�d��lS�;j,K�ʴ+bZI$��>�3�p������]�����9;۫�ù$�`z�k���O?<[c͐S�1���<MQ�}gH�Np��m�/��CV-�ח��?U6��,����Zx�縿��F�uk1� �\>�u$l*e���pC�=�=�2|tv�e��7zn�;�L:�g�2��S޻�``��V�WNY��$ޘ���V����j��(���6d%�ك��:I`kx�EL�ڸ/ȈF�������X�gF�KU�1��SE�t��z��b�bg39T^9����&&����G"� =�xc-d�2qrz�ӳ�[GG�}~��ȭPU��7�T�䅒q����bJ��8�?�in�C�W�p����u�,�/"���g0D�
�2�9�D�b�~R6�#L- |7�����c�Ym�l8h���x�tm�*QL_�M�u�M�)["����VIwğ����N슓�b����&��'�)p�ld���Nd�J�^������#�Y��<��7���
6�+G_0g��t�I4	g�홁F�'#�2�2T:Л�k���G��v#!Zd�+Χ�_Ґ �oc[�GМ'��g��_���z$��E��L�F��`��i�.�!�c��%����g�O0���k��f<�b�\��X�ڗϸ�)�I��BE���Ō�(%��й���7-�Qv�]��M7;��Bަ���{�"�$-��&�}���˫+y����$<�:%_��
�zξt�:��<��,5~Y�����+3>��1�J$T�6 ���m¨�>�J&x��y@Ȥq�haQڎR}��я�;��{�g�������"�i7B����`O���z��mp��TKl#��vO9)�ʿQ�w2�#ya"wC����D�
TI
pQ>x���-XV�=��!��x��R��j/�H,�U=�2B�e��v]n���K9�yrLƠ0�9�E`q�Pǿ����AZn&KX;��?��˦3�?��\�5R[�OeMe���øH4��/�=@1ܚ X�,�y�]�~�5�T����2!qG�xx	v$���ڒ_z2���^ϰ�=���v�Xۓ�����R�Z�e#�*͊���*�����w�>��(DpBB@y���g�3�Y��^�t�X0���)7W��v;�%���e��h�BIr=�����KH�$��_�݉.��ˈ�������O-{R~��y��5Et�푗lG�K���o?��-ɀDd�Łl�]� ��	�l���X7��5����jZ*�N�GϤ�9�/O7ς��P\ݿ: .[�����Bq	D�d�`x����u�������p	v��"�?g[�͇�3YHh&���ښ��P�:,8����*��$���OD�g�Y�|������r�NBU���޿����(�rC��{���S)�ܝ��l�����C��Ś��i��zk*�<C/�&��$�z�r�Th��E��W>��V^�r�;z+�޷h��`� �%L�ZL���|�ߡI�B++�Y���Վ�,BwJ���x`���XI��c��0a6};#�Ժ�)��Xt��'��9��c =S�{1׷8��m�@)����X�i��c� /���)*�n��ZM{�Wd�iI{\6¡�n�����@�=3G2S�A��_O?�ș�O�s�f��".�K�]�Kٴ�R����)<�~�VK��.�U�h?ݾ��j"��%���â��YV.��j �%��d�����Z2��'f-�7�� ;�/��RRd۽�+`_�d�"��O_��A۵�]��|��e:̂�f�sᴚ�
���&8LϠu��+��ו�����[��`"�����U�p��-v����Т]����۫�0��ţ�K��\$��L8x�o?xeY靟I���H�-y��1�7���ˏy0����X�,�[cC#��O������*Y�^�V�L��I[�J�d���i�vEl	�)k>3���f]K_7���Ȳ&d�1��� ����=��\؋\���|���$�y���K����4Ǣ�x�B�:�G�z�A��A���H�������>�Wf���*d&����}�z�杯���q|2���d�-IWQ�vU������W�b��J�,`S�*Yf�d��M7�h#�y�6�/��J[e։i�9</�1*9��*)ED��H(���P�UBa��VTUT��{��n8���ԘIQk��&���VC�O��;���߲� ���RNFI��FLm���0����jw�{����*���5X������(��^�i6�d-v)	���Ӧ���e���2�r��$)|�����5�_�q �4�hZJ��u��.f�&}��"O��m�
�� k�`u���T����F�"YcJ;�&_v�I/u?CTs�Y2Ӹ�㾬�q/˅p�`��Z@eD���Z��.���/a
w�*�n"�d�}���"Ms�9�kk��L��2'r�M殕���#�ᇶ�t�?F�g���)eU���*!��3,��cL����X	KY��!Іs�*������C����֔��Ѽ¶��5�s�%��T�"ՙdZ�oq(C�c�y��X,�壙7h��<x�WJx��R��MyY�+^��Y,��H!�����S1u\(�4*o�t�f�Z�	K�[ˌn����L�Y���Ng?����"����5"M�x��%9�8�N�����I���gZj�f6R�tE��f΅~e�y���	L!qЕA�r,��㫘�2�Ҷ(H!G�y�����E�VzlQL�i��?=�g�66���HJ9X-��d�+���Q&,����|��&H�����(&3�5��df�ݷI�%Ϭ��bA{�ï�^�)\�S�=��3����ѪI�hH�e����凿�*`Y#��'�:�\�R�u��N%=Ѿ.��W�0�L	T���D��P%m(��N�C�(0����s)=b�7$*)��g�c+�^�v
��Bh6�����$�?����X�s�p��ꪓ�r�cś�k�tշ�������gi�A��/ro&6Ȣ�����j��;�[�����`mx��1[�b��D�B�����-��&V�S�G�{��
9$�#J���?.5��w\8֮H�^.��m�%�)�,+c>���W�kf�f�m�3��4�R9y=(�y1%����m�y��k:-R���2�]Q���l[�*�*�r�T�Ϻ(�����ܠ>GP�K`���O�|
w9��E�ў��*�E�M�����US��fT���o�0�rm	l��jzR^F3���c�����_I��B�]���5G�4�Rpq��|�.y-�#�h!��ṳ7���Lf�k�p�ρ;�+b�������������8D���ڕ2{��e��ۓ�x���:�mֿ�"!�� ��1����mc�,��;|�Rd}N�)+��C	>$	3�t�|��MD�̶�]��Ă��"�`;Sf;R�u��%��<��cm|a����x�	aݮ'a���9&�SJyf�ڪ��ʯ��q ��4�k��}ה��x5;���r�U�}��1�h�Lx|���H+Jt���h��w6��AH������s�|4}w`�h����|v�q,��hY�q�P{2�HYe&w��~9U�0�L64 �Y��/@�؄���S�"���H��j����"ԉ?��vIw�Oj�!��9��,�M֣�\�\ץ3�m�kb���)R4��Nd�z�Y�Wju����5)��C��m�8{Cw�5�xSl�r
_3�KP��D���qH���XƆًu�q�¥fQǕ$�����������t���g,���^���/O��}�`u=$nb?&�V��<���WnG*�vW�mMCav^6H�*�ƒ��%��C��k���=�\�@��Bs�eQ����V��9x�#Yٟ��m��9�DHPv_m��߱N��51�'�,��CP���$�>��C����Ur���ݎ]���Ӷ��K��[�:q�:}UA!�Θ��h,����'7��4se�I/d��x.!��[��#�SR���l�rGR6�:���_��⼒nt�3-�-��z�'(2���5�O�獏��h_]�^!��*�1�������:�����;�sn#��/$v7���2�Q��h͛��}�du�����WY��w�p���	j�nB����-�ȵ���?謨��G��bn��i�-U��o���إ�iK�Gj�{	�4TD�1X�w6`2T��1'tO��Vx�ȘZ����1ĺ�L?�1,���
��鳷WN?��t������R�+,IYZ6�� %ˡ�ǾPj�v�:�Ǚ.sd���~W��pޤ��g��I��g���J�u,�!a�qB��I����l%�8G��{�����.��k*��$n4�7'�V\�M��B�P���2P�
�=�S��֧@*띘�޻���-��$��.O��ץ<�;��VUS�	����3��"�Pg������5�^r`���F��y�����>牣��4:��]�Y�Y���S�\롪��I��"U��F!攴6�9,��T�����0�����{J}NO!�'c7O��f�Ի\Q^��Ԉ%K���{��6�?�~f�wR8U��xv��1�s1��H*�[6T�H��B�Ew�A��㐳�������i`�>��3f��%�ȁ�;L�wM>����������l�k�����2��"�Z�𿑑TW��PK   WL� �� �� /   images/3344f319-942e-4277-a6d0-796a8e5017f8.png��S\O���]���[�H���n�4��.�$��>� �{p�ep{���w����~8�u��սW�����O�X����޽��������T��������S[Y�p����;�wd?L�;�3)�<��y7��Y����lh�Em�⮬.��r�-�-pqĊs�r$%ᆷ������r��9c��z���pr��������.�}
g�:����#���mx�Blx�'������~V����������1�����%�L�(��	��>m!b����������0������f�0�e��>N�#�/�ch(>_���7�[��῵d�p?�������߂Xd�,�K�c�{�N�����U���k���A�G�*v���BD���Rߦ����Y�z��������?�����W���6 Z7C�����T��E)��#��mǛ�����\�����F��C�m�gX&ο��3�l8��y� �����5�B�r���������;P9�1����fܒ���о�cd����@��s~�*�O^m����O�

zn�x�,W>�cc�NV��Z4�_����#���[�әSx�c0͖>���Dّ���O�e�I�x�HorE��q�$~���&ۀ?k����ổ��rC�k,0@"��撎W�]|�����*�Q���9���p��뎞��>�쏷��X�R��+��r�cVW	x�#~�V��L��x~G�n��_z_ל�V�(�O��%j��潍1�����!�F��W�,5�����#���������r�D��&pA0��5w��\á�I��8��4��T��A]�̫�˵\&�|8�h#�߽�Q��_�Gc7b@A<JBNf
�x��?'�򲳳֗�c�qQ�� F��#Ɲ��Ӌ�;.lI|����`��D=U����퉏��d��ĵ6��<�쫰�������1vb*e��ҡ�ɸX��ᤈ�X�<Oxz�-Y�i3E�)i�'�q�W��_fiS�&�5�K��|��LL���
��AKKK�_�gnr^��2n+4lv���tZV20 �����%�)|��D�r[?S��FJ�4@O�TTW��h��d��.�������ٶϔi�mg�1�x���b���Ɏ��E
��s_q�r*c��g�L�A}��oH���@�HԅO8��I��p}Q-'��thLJ�;">�I��O0:�"�m�����.�=Ϗt��f ��TJ�X��>�9�˅��$��E��x�G%�Y!L/�Y�u��OfF�O�:�V��L��4��К���xzm3f4~����w��H?��7���H�i�BX" ��Q�1
�1�٪���<�m�E�������W�m��ȅ~j:W�����."F����&�!�W~�N�M4�ս-�v9mgG�)g8�װ��[��S�	�;�e�h��Fci��*5��6�pF}�I����GQ�ZT����bޤ$k׼�h��n������O,By��d>M|5�Z����U},��B�F4�%fMaR�:�ò�	���^-m��#�$��uVO���4��L�H��iu�~fJ1�M�w_�k�,���	L@�c�)!���A���6 ;�ev���x�ޭ�Wu�Ȏǁ����HI��(�~YW$M-�H�Y�G�1G���zg���jY�i�d��LT�:s|�w���v�8�:�������F�'{�kx ��¢�H�p��MK�%u�Pu�R�̾+�`2F�Y�$mm;c�Pˢ�72�����OYl���8�::8`~ћ;��+ѫ6�_tZrvvV�d�m�r|� C�##�YV��3&��b~- %p�,\h�2���F����M��N3���<[��`S��ںUGG��<wq(Z��l}OX<�V�)���Sf�!���\�U����3�H]���}�ڽ�&!�������mZ
�4`��Q�5�C�
�ء4��F��L�g�x�� !l:1�e�~�據��w�7����.�$������;�d�������A�g�/$��mQFʕ���q��KA�NBI���1珁�y7t� ���#�`��OR�i�,N#M�Y�Xƾ�Ԓ�qj�c�T����C�S���}YǗx�אӒ����\�E�w�5���,m!Q��	����'G.]��l�'=<�{�0�Ī�R�#��	�%z�2Y��5�K���r�`�*��X�?����en
��9:"0+�E<���Ë�D����q��2���FG/�6V�\���V��?���1?�?���wUPd�0�Ǣ�])�2�4U��tv��g-��
�,����D���%*�sD�A81r�}c�K3��IA��PH�u#��%�����nc�+���($@�@���n1���kZs�!* �[8:£w��u��|X��[S:�y��W�hp'�({8W�q�د� �����.�0��z���:���н�������7�yo�����0^������'	��Io�?�?Ʊ�gp�IO?�OR+�2�ST�̆(�=����~�M>��P(�`�Lg1�U�>��Y�.]�r--/�z��}������N@"~:���966f�xs�LRUU5�G�LEEu)�	�x��ubw���D�&n�^���۾>|�/P�ԡw@��������r���{ߦ��M�i���G!���Aq짢#Ӳ	�y5������=l��^RL�ԏE_�x]�[�
�=&��Q|�S
�?�j.�9z�ٕ��j�1$������pcJlT��tں�^bc���ۂ�xV��v��mhˍ�K\��`�a�X
�=u=&�ט\�w�W��
F8pRH+;��&mc�Z,�xQA��a~�i��׀y`�2���Ã���!5HƧ	� ay���xR�K����7͌�[�|�|����s&bI�h�!�0�]w~E�1_�!�ժa�nm��&)f���n�!"�y��Ȱ�3H��Q��A���Ӹz_����r��A��Y��>7�t9E����@�~�w�|�2��9���!�A�w�g���0tw[�5�0�~�Z�)j�t�i7��
3�O��y��K�����������5�9��p�,��f-������#�30F_��i��·�3L~s�{Gf'b�g4';�9ă~+�}va��d����;��Iy����X�z�Qp�9{Xj��j1�3�6�Y�9��P��ّ��H7��-�/�(��U��2�%})�r�7Q�����ެ�I��� ������Dk��%)"+�����%u�7�P"�~��}�h�d�G�.����di$o��#�b��1��C�OE���S���l�࢐A}������/�Ce����|<��\u�_�x5�ph�L:�ceuLL�������s*�O��V�ĝ�V,�qx�F?���6�z�2Bf���g�բ���1��P����gd��"V���
f!�8�t9=luK���+$0�v����7�|PPGn���=�_B��B��a[`F*ϲL��i��YB���Ŷ����K�e����� ��Eb���E&!�F!!<���`��1 (XT�:�^#<e=�d"�agn�h�R(���1ch�Uz�D�gJ��e]3</WZL�sR��%���v���g�;隋{���x���.S5,�#cCmؔ�E	�)�dG�D92}ţg�?�b7�\I�(eh�{No=D1�g0�]��9$<aF<�x���̜�Xک0��P!3�E��2BY��
��Z���'H�|"��6�4�6��Cw�����^K��hn�E>P��[�]
� =2���(����I���M��b ���dT�&�Ў��ȸ�G�Ҳ��J@����lF�C�_�I�Ƭן4�Վv����wȘ����[n}м��"��q�q����ͫG1�զ]&9��.t@��K_�Q�֛3w�m���&�p.B�H'C�%��7�����<����v�kM06
����suR��R�H��C^��,����$t���DN�/i)�X�=�S}/f��I~�eGS�db����"ʷ�/�T�#
s�sr�L�<��"�M�&��U��g���|��-���y,Y��l�BEd0�`���X�-Ӧ��!��zjo�˹^�$���ˏ�Ǯ���R��3�ȁ��+ԑ�mR�8����W�o��4{�W�B��"R�Yӹf�mU��}c>�˝C�^Y/���k-��)�l�>5^�)q�������h�f�gڣ?�s���U�}���˹�9
��o8Q6f
�J��%��0*�������[�\���v��!1��*CIrr�ª*�D�����f�v�F5���"�On���zy��� �i�;����yB�i+��{�wD�.jI��Q���~S�T��XxR��ɩ)&jLf��C>�n���W���y�~�� ��׏���1�
��inal�=��؆݆�gl>]M�7�C�vG'��}�7{~h�u��}�h�S{�* i�@����2[��;����N+-d�>h��6ĝO��uu-'���]��Gؓ?��*�܌�NV������������o9(3<8�6?���}c���D�΄�\ʅ��?�@��3���\�!s��D�Ł��]�?�S��J�yk�_�&����#6�:��:���>���R��p)7&�=�v@��xօ D�X&Jw=��Y=鼻O�c'��`2m^��X�RwZ]�!���Sn�c��n6���W��p��{�s�N���T �-��Zd�HF~W���z�9_�WA��s#����K��ʖ�~V�9�'O���s�?4��-r�������۫�q��Ʉ����w�>��؛�=��j��>pa�.#��p���
.a���d��3���=8��ǋ/Ţ���+&��Fa�!e"���G�~G;;;\ˤW��x/5@g���K~��A�{�N�&U�g�o�p�H�Jz.�,
?G���0B�Eܞd��d1w��H�):d��SD��6l������o�?m%�M�}"	�G{p��`��mMM�	OtϐKX�)g�/ ��=�|1�3���\!k����F$봴�]8c�_|,w'a�g��\�sb/nJ�TY`�RC�fHm��CQ��H�N�Ф��b��,!ی�]�0�'-Vb>�
�*��F�6�u(�D� �f��e�.":��9ʝ������P� �_��{��i��M��W��T��&��4�Դ4�pm$*���d��
�n^�1v���Qy��IM�,^��3%V*��}|�R;��slvq]�f� m�~�����{߻��a*w��Ӛ��$SR�L�J�,��m?w�x�P��EM�I1���-;��ˢ���(䵓��i�:��/l��L�G(��)S7��<xy<�^OJ��Amʻ8g`�Y��ћ�grk�o3h+��6���ة��KְU���������5���0�ÄBh"b��0�h�3�U��?$	�`��[t�z�㷁`u��w��[%���q��E`dh��kwvc�d#�����#';�M��R��p��Iӳ,0;]���������[[U~mT��w�C�� ^"���\7e�v���^�ޮo%G�(�A����l�n�W�An����wbs�b�|�HR���H���Xs��/��ެ�8�	Q�ф{7�Ɵ��^��u
�b�)|<��N����-4USZ�9�kк������!����9.N�6� a�
�~}�z�ો�	钶���r
E�ӅvjRTz�A�㒷F�단
��C3;Q��Ev>��p$��Y��ܵVk��HY���^W�+ji����:�阖\�b���
�,.۵�P�Vdt>�1��o���,z�ȕ+�P�K.}�R��$;�fg����xP'p��'V!Ǜ:�WAB�#��g�'	��$����@�E�Q��j��G�H?��M(��J�@n�\��:��Ojl�
�A��p�7����F�.|_���-�2u�ʡXq�\!^�}�һWS�G���+�c��K�ş_tႫs�o����Hkϻ�W�Yct�U2y�F#{��l<i
�}	'����(�O��G����韅���..{�>��Jg���H�g+��_�E�ز?eD\8����.���նgk]�m�.ܭ��t��8w�2��A�I�+��G"z�����ޣ�0ˮ�58���2�5>p�?T�l�ɐ
.�=�(*�>0BE|��Z.ʎv|w�Y��ų?��F����ݺܱ��Z%n~��SD�
�C5n� �mK��)>G��%v%�\���]%�,�,���X>-�a��O�f�ƼG�fw��d��9 >3�O�\�c�/Ù������a��z��=c�"` ��zcD\�@�T4(��;���M5���<�$�lUK��i��9�T���S7W>
�g���w4O\�	���b���3Kԓ���+��v�5�P6���r��~�j0&yK�L��~"d 
��ы��l9�C���ۂ��3��pJ˓�ƭ�G�6/V���~9&�3�(.�UFSM����R�Iy���狶C�D��D�`�s��!�A�I����P�� ���v��%��O��Y�-1�6��]t�T����^�&�2A�t���G��-�F|Gw�v�%J"i@�%�$51�:�ƜK;:#7�3�\f�!�ǻH�ݥ�YZ��t���g��Ҷi���PX	2B�J&b��<i^'�V�<�
Xbfs�'�0���J�/�geN��q�$�~���4w���t������}�r_��]���>��0�s�J���/����y�0Σ�M�ҥe\��}�y$�x$ψX���������wP��[X@��Q�XQ�W{����(���gU_?b�X�9`:)q	7[��MV��<�A�m��-���QJ��|),��TW��sa��ZA��ѐ��v.�����@#8?`. �����"	#��N)�Jp��C�&��=��@�u8��d�ڨ��R�̃���f�	���&eE?[��N�w&����u�h�C_y�#uuq%%�+y�dۈ=����4�F-+��I�T���hZ�1�ȭ�R�Ҕ���N�٬6�]�zD��>�B�=B�7��e��gۋ��{�'���]S���΋{�!����(��~�e�9���LP>���u�0���A�5�]��R&�Ad���a�J,�J���bh5	�ݟ���6/͟��P΂�Dh����r��"fC��=�zK���~�%u,��������?4�A-3�e��,a��?�yN�B%.\��x�0��/rә�^�Ri��vVݸ��"R'���k���+A ���	��=	+Bŧ��b�7�DB��������?p} ��7�m�xp]E6�;Y�kPH�94�W!K�����`�5�6�;�R��BH]ڠ�NK ]�)׮���②�t$������v�͛�吱M������8R���i��d���xV|�<�`���K����ꮗ��æA���a"��L�7#E��?p$>I�W ���k�Q���k��^�<+�w�)�J��G�E��eͬB�Z�6�(��6=(w��5�Yn�!�&�:@.	$����Ձ�ȨՏo�;�cD䂯�������^Ϸ~�i����<|�Ȼ'Hr��v�p�����b�/?�PO'��Yc�J-] {0��J�W����O%���]7�V-��ș���Νߐ^�k׳��¨�ĸ�QLe�9]�A�aҐ�Y?��s�*WO���Gz��Q`�Z����8rzМꃥ2%QPT����B��+%����)X3��6��k�g�[�C�Z:Խ������}8��q��`zMr�8������i����1ŏ�7�y���B
qcd�,��\ftm�9�~a�	9k�4R���@���$R�ն1�KXu[U:	ϗ#!���I�j~~�1՚�- �H����2u*I]��-p3	R������Q���Pl��,��b��N�9Y757�-#����a����|%;n����M�l���A�̽"��+�G0$J���u��U�g�Λ�HR�I$γʞ`u5u%Y^����(��3�Q\�?�����$�/k3�p�iI�f)J_*�,5U���ߘ�X���߼1��,�f޳���k���ɐ�j���HW�����MslΩP�d�S�3���U�$�M.&��Um.�֗���Jʎ9O'?g�CǇպ4=����#un�+�������S�)Ƈ�>��Q�c$nz� �oW�1B7�cw\���L�6�{�N��Ki��`�[������  14��3@r�;�er �4CtE���Y��i�y�ɷO��Aw�����*�=�Բ��{�#�#���(� J�rl��7�ٽ-�ֿ��-v�CLg:���C7�^��\��M:CF5+�$y[�A"!(�����t`����S8���q@�w��n�����߆v��P��I����a8�etbňT"f��:�џj�<�+
j�p��hH f�n{N&��Я�����Z�{��-�~��◹��eo	9̒�rK�<�,k�<�L�^��N�5*}y���_'���!��;N�m�۩��=e�۷���96�4�HD{����,�J�ϰL_��������C蝠jRQɷo�c�u�d�5��b��6ʌ-+j	�����G���lҗesx�Q-_ mB򶲔8�B�ßӥ���Q��u��ʫ������~�Ի��q�~\���@��B��:���Gz��c,͞Tk�|����F��n�k.��ٲ�e'=��i�M�ئ<� j;��u �����	�?l���\�=s�F��9����j���&�I ���pZoëM��<^&���c3	�W|	�k�Al��^:d8� ���ԗ�P��?�U@H������n&�t�r��,�B1��|���N�)��|Eu'���q�����f4�5� ���<eҋ�3��%�~~NCݿO�c5H��B�SN���^�4�a���8�oy���g�qO�##qBA�}S$�a�e���Y��(�$�����Jۨ��p����F<�EQ�����4��
a������ԁk4���r�I�K��I���O�=�5��:B�z-i}K]�)�Q�����d�^8�ڈ�=�t@���W��NXF��C��:0�A�h��|��)uoDO�f��X��6g_t[=��:V��B�q����!1�����3X��h^��2.��&���O�^�y��[�Q��ꏥ�h�(=vOm-K��u-�t&i��of���nD�SO�Sqxjm*�p�6�\�%��E��J$_�m��X������O��t��pR/��9H窄�z&g�qxs3'�f���(�E�d�Yk�d3�t�k.Q�XS��9͌q�DD��=T)�ܗ4v\889���zP庑�mz��P���f�H�{�
ZB8�U��T-?NبQ-c�N<y(���������g�!�G��P����az�ʾw��J��=�vە��ҝ{�Q�O��ds�E�
f��<j0�j��v��^����%�"*f<�enA�lv��X�t��<�/k���E��o� �op���6
M�놑�e�dE��2%@��,��M����D�^í,
x�)�|;�mB^������8��((�����w<�$�������V��q�y�)Y��`?�|�S	�f$	���1=�0������W8;��Ok�q��sSi�Gjd��C^�G��?�yprU@UÓM���A%�C�Oɞ�f����~�S��DWy�8S��9УE�wjŬ�anI_��P�^k�I��?�Y�s�� �~��y�ȟ�w���ch�-a��\ �6���L�����*�[��$�b�׌��v��e߱�#!W��Bɤ���ل�^8��F���tbV���s
��P�/ݝ�T����[8�U�,8m��!<x|k���8����Ԓ[��8��_��3�Җ�}���e;WWy������~-e��x��^o|�uu�D���9!%t�SF��̞�:���8R������1I��|�r��{ܙ)c���W��	�&W�ś����tD^�cy=����3~+M���E�;(�CS���1��ub�U�-�-��d��2�7U�!J����H�nU��˟8�ݙ�:q�6i;H�Y�D8V�"w�_'=^�(��r5jGNtڐG���NPW�0BP��NIE�wH�ʕ5���32�@�L��f"��uO�Ǿ?Ŗ�%�5I����zΓ����ww��x�Hɵ[-�ge�A����W�!н��W���򄡉���
��w�TD_�]��+7h<U�/77�S�|\8p5��\��9��]sXͷ�Ǆ����
Y���n��j�'T��6���a�꿯D�_/�Z\�}��e&?��/�`�g�uu��K��t�4:�,�O�
Mf{�!hsr;�:i�ذ���O~�C I� �pLA����Sԉ=�\4^��^��@��(nT��=֕�S10�Z)	*F��q��(la��*W��$4D�%hP�˾�Q�U:�ܼ<<l������q�ξ\��J��u4:��7�O�l�[q���;I!��s���Ui������f~�W����̂ʒή�	I�"�nV��C���Z���}�����|{�ew��:`5�:%�V�m�pT��X:�ĕ���SW�.�Gg�����-�I� �Ư���b���]�Cx��1B�oq��e� B�,�y�'�i���n��@�3�']�z�j1f1bBɻ����-t����}g�t+[K7Ms������yl�0�����~ߐ����J�#�1�a�4���i0/A@��H���vT�>�R̘/[Y����*�A������(<�|�Wz�~6�[e8YaK3T��Tŗr�������7�������OY�0ir\[%ĉ3�۞��k��J�����t�;Cj�����DG�r+,%�	K1�X��3��70։�TQ�F7n�����P�]�X�a`������!�+�f�:�9��}�:�/���:��E�3��^3��l��/�I�,�sT-��D ӄ��|�o*�����l�9�y�w���ׂT�R?�Oz4��#����/�w_��v͟�� F��c�c;�[��-H�|7Ц���M��r����w����>��Y�#��,����d��'M�g5/����������0�e2nm����lq���}�u����R�J���6��Z���7:L$�r�0o�:)w�ؙe]��CDe�=��xV�qe��&y�����%s�l����t}4Ye˝xxpwy���ٗv�LYG�?�>�L�8;���t��^WTW�V�,w��֖�?���=i�=���=}Ղw*�M�q���t��6	`µ�������;E��!�R6��ʎ�	}׃�[}��ɎW:����Z��݂~[�W���Y�
�n�wD��ǪW��& ��q��Ku��lu�<J���"�O����PB�N��>�������y�Ϊ��l���Zҁ��e^�^����.��4�\��G<pu��o�zj>C��I�Q�M�9q��7^�#����#��J�����W���}B��9�t]�U��j>k�<<'��C3�Rg�O"?�nF	<�:ܮ����ޫ�$�?\��9��0��s�f)�\�g�:�A^��������b푦T�ti�H���@��ڌs���p툡^=�8��S),�o�|��/H�?�wX�����Ώ�&��]��g6\���ƫ.S�^b���=�P��.7!>�r���prZ6�O��1�m�Q}3�;�Y�tu��?)4��Łe��	)Ivt�.B�|��k�]ʵ�j={~y�d�f�5�RewW� t14�,O����s�D1䐠k�'h��T�����J|�U;�1��/͛�*���<�+���kg���c�o�P�M~k�̮���T�#�ϰ��1Ϳ�+Mj1ǽ%G���>���J�]Di^u��ln�<(3t(F¸�(/��9����y0��1�d���QES�!�v�:-�!=�2z���떫RI�`��XTSyU�B��2K�b6���H�z��]��N�VB�Ό�Z�r�fi��u�ksz������cQ�㐍`��}F�W��쬗�̩�Z����,�v��֡�πK��homm.�>Z��4G�x��8����j�F�y�6��t=�]�u蒷�r��LR���k\礥5��[ ॕdrn�����Ԡ�ڄM0+�.SV�3��EfeJ���y&��
q��e'A\�D�@?W��!�D�o���k-vXkH�������ʘ�c�o�ч70�=
�b��&ja����r!?� 4����3�-B:`���bv,��&��\�"N�ə¾�پ������N�t?���M�MF%������H�����k���
漠�����!��7���ja�$p�)�g;E�|td��+��-�(r��D�;[b*�6ySiH42A$�\��z�4���?B� �ti[B�&[��ݎx��2���7��b��yVz�x�`�h�h���R(O���tmX�O�EV� `�kt�D�Ҥ��Q�WAJ����k�A�j�'����v'�=M���x��{T��M���'��א�D�B��#A�����se�����|(�%��$�r��R'�]!��W�Ю�]v�.��=fv��������H<���y�ʥdM�+F��_��B���0=JHd�lx�<�#��Cm���=�飼�O��No����s�I:j�c�,v��z�	�y���J�@���+P9�ӳ��D�C~�zq6�lk�D�����@�����@KZ0(1��9鞽�")\�>�#�f�:��Ye�Ƅ/'���e9����0W�l9�Ş1GMp�%_�N����LCG����p�G���0Br�7U�»\FF�c�\J|vj����Ƅ����?aӭ��ӈ�ۭ������f��l.DN��'?J���$���uᰧs���=/y�c �A0�3P�`���!s�P���D��o��^n�p����`n%�[IF�^Tt��5(���궇K_�����w�T�D%��;zFt9��u��]��
BnȤ�a3��(��^1cݺ��(��y��K�à�������Ce�-�Y�E�{��I��Y�&�md�t8���Ku���p�����z��2b�3����Y��6�#���N
��S��gW�g�������_vw�_6�y�#>��5���A�f��I���1��?���#�Ǽ��sՆL�mԭ��o�%f��U��{�.�,�̛���_�q��`��#�~��d���bT6����!F۬.��UGF>%,xk��q��C�O�@;W�:`o���Դ5Y��<�o[,	y�A⺯�c����.yȔ즜�d�+)�j$���g8 0YHww��k�EC�q4�����{�Iqq/-��$l˗t��B��ϐ����^����bN
�������gE�׃���g[�~��cW��~���{,�1��=�%V��0����P�׷�ԐGn�������VRv=�R���pj��y7�9}�xq�`�Z���r�ܵ�ޓYn
7���b�����?�l�#㮣�(jTY����6p��F}�c��Q1�3�g�j{�����'�����y�i�r}iBVN��>z�^⩊TV�Ψ�^t�W.���E�Sd u��.�3�1f�q�f�,�g������m����+�>*Q��&�+���X��x!a� $�C�,\؆��N�A<!/@(�H��^jǟ;t�w�'y��Z���A���A�C ����%t�w�.�_��S��e��]گ|��>�lvY��.�Gה�'L�0��w�\��ȱ�����!���wo�!A�nW��)w��`�`ũ��?��r�1urF���y]9H��8��W�ie���n�f�pt�ߙ��Y��r���6E��5�8�:�u�}z���;���j´�^��<KP��F�8c��$�<�wG�⣩��cUn���
\�H�E��Ռh+ж XIv֙)+�l���x7SP 8��%� �uԫ�b���$ߐ�ϛ�P�t<e��6c�H��3	��z]X�����b�J rJ� ����{ yN�/��"T�f~�����9i�9tl1������ ���1�EZX��Xr^��or����H�E��׉��~�`���4n0�����0~|\����gx�8B9C,���ړ40|)�e�:Q��W�}J�EKI"�:��}v����S�i���
o,/�"�h�#�\@%�R��@{�5��)��%��C�xuzR���%���B�x�Rw�Ƹ/OO}r��f7KP�z&e��!1H~0´x)0?��~��"��?�������������|������ka`�8��6����b�B%RXP��M���Ay	���b!�����j����}V����MN�T�X��	�|>_�4jC�_�M���͎�G���Ǖ֥�y�(A7��S���&8@�nByA� �+�?�p��l�v�����w�,��"&��}@?�2Բ��+c�s��<?�f7�8�����@�Y��;s�@_؉=��zQ*2�V�O�2��؉+I����`i#��p��ˎL|��m�s��C��}�h��qm���5��q��Tvg�zy��v��V��sW�QA畿�+�Z�.Y-q�CqQ>p�c@(B!$a~��)aw`�Y���B��c�Hg�:�{3���d�i��Qo�u3����~l�+1�Wϵ���3�T�a�EJ<;��������)���F,51���u�m�e�!r���"pLeݮ*��gde� b���v+�	�����Ĵu��zVt�K~)���`�Y���q (g]��X2��l�#+C}�8멚m��x�,5Q�i�Ə�Q��I��f��[�q,�b
�W��~�Ęb�%��ހ�N.$���$�Cqz/��'Cd�+���}����*afH�\�!��� �KZ��C��>j��Bn3������@Q�%�u��\�����*�&���[��i� ݭAy�� 뾑���4V����]�A.�(:���!e?�ۧΓ�G��`�O�)�ܽ)1n��GL4Q}��D�&�t4�I��	�6/c0�t��L���	�Q�7�݂{�d������u�(���ݒ�9��͒},�ӐOQ���t>��Ԗ`��аj�vR<�3-z�I����n�ĤoX��'H׿�P%?5_�6u/��eE}�f&A�x5 ��~�y!����r*i���5�ʷ�Gd���J�;�j���?�%�9��ft�6����kJ�a?�v=�o�	�z��*C��@f�ZrE�`�"BS	S��;+eG���� ���c�d��������Lue�!�L�Yv����Mв��T��Qп/)K�P9�������F��ׂ�����m��_�PGc#YUi��`����G�������y��s�ʠ}o�mޯ�+�i�C��5���0נ[�vc�x�Ώ^��`:p���T7~2F�%�gR���@N�ۄz����3���<�A��2�	v~���F��7G�����h�&�O.�Y�ƽ�e#�l9�H�O�	7nN� R]`/��	�g�g�ɾc�aUd[,�$+:
1�;&���;G �UU9�x,ň�ĩ������:#n���tK6��UW�� ��b@���O���A�h�@vMA��M� >��m���fW��Z�)����}Ͻ`�������� =����G���tiMV�]��^���sCۿ<���y���~���@ƪ�|~�~7���bX�$���R���h �P���9^?��o�N2��Z��\�x}
Gq�������I/T��SIyhj�J3��Z�zL �w^n6��reu���P�e��-j�_����f̤�N�$I�_u�♇��c�s"yCJ�e��r��Jz�Ih�>Q�ϩYy���2�|
$E�loq�r�n���$^ψv�!��O������6�'`�7�8���1��MBX�<��7�u�$.��(#�tT�)��N���]��-pu*k
%N��Lh��C/�����K�]�i5$�є:�J�wҕc=��3^D�v�H���2�>FJxn�Սf�7S��[�[����2bqGUĞ/9��z/җ�	�x�:C� �uC���K�+�ŝ�k�ĜO���&��(�x2&�J�-k�?�>L�7��7;��[�zUT�S��>�^MMΆ��ʄ9&��[7�*�-bD�2���%oc����"wܜP��_W}�c.f�8_
�p�$��[���\.F�	3ڧ̬M���8��i˪�[��vv}Uͫ���5�vnYLʹ���Y9��B�g��:n&�`kAG�O��惓p�X˖��nO �/��֛i�`�K3br��:��2��]�Gh[[�_9��}*�D�����s��.@ѿ]����|��+�x��J��4o�Ȋ,�t�T��ĭhoj�,��¨���]���f��y�AlغY�R]�p�W��#��� ���C����?�'<e�M���ۿ<��F �G�[��]t��v
���J�3ca������!�s�54!��о_vKڱe��v��v&ο�v�k��-�A(��-Z�S�,yx�~X?\o f��\^_px~ ���l��@G:#K��0���@���o�����
���̫�={��.��ek�VX�N�|��q�R8���bݺ�Uvͪ,���ի�Мt��U��N�D<����ӝ���@�]��K���\�l9��ۥj7-��ef~@&t�Nǜ%��i�݂n�ch��DPSF"�0��hY9��*�X��׊l]sP]U����5�)U�����0�p��$�N��>y�C��)aYN�ŝ��{X�Gc��C7EQ&/~V���/a�_�)�L�i]���/Nƌ|p�->P���J�ֳ��qP��F��'Ǳ=|�\|�4���"V؛��/>�����d{�d��n�b�5�;��<t�_�>"����6��Q�09���6�9��0��{��S[M'�x�ϟ�og�D����(7��A�b5����eil�%�+I�@ǩ'��w�yW
�XƐ;�,[�B����*wVѳOؿ�'���������+�#�k�E���a�j�!;�h�l�����Ǟ��۶�����R������36��*���Os3h�������.�7�~'k�i�s�櫹Q��������'��ش[���/��o�.��4;F&���7���MW���L�9��vy�	t��.�u�޽���������d%��s�Y�(<����x�7лG7�!���e����Ceu]a��|y;�א\z<ށSO9Iji}�UT#����O�������[r)������y�#mf�m/��V�]m��&ᾫ���&cҸ�X�p~\��`�H�]z�xn��,\���Ǝ�f��Z�9驌�JӃ��=�M���#T�h5ĳ���<�Q�pQ��j|lRFC*��
"oE���]�8�<�d<�Q=`$f/]&�ĳ��k|�צ>�x�p�8��k�$O���P[a"�M5\-	9��@Yda����+!|V3����:׷S�Nf0�Ƌ��꦳��v�I'�����]W~�`�=�qL���EϮe"�eQ�_�R���i4�h�b+.w�cc��ȤW��ѷW#��G�qp2�TUVvE�~�$5���oHX�[�z�XIχ�0��s�~>B2k�7O���uS���ؿ<�JG>�D��#�/l=�K FF0��-m��8\��'�+n�!��rp��>ڿ>�R��{�(�������>����d&B1 !Hq�R\��K(��h�����B���Mq����s�9[����9��_?��]�.�o1ke�d��s�<{��j5��RQ�D���Qͭf#Z�����i�8#��]Ώ����ZP��l�*1y��\�I�����@��HD�0�*L�g�\��t	�B��i��Li�b�r]M�X>cM�X��(Ic��뛼�lܧ�	�O^_^�f-���J+^���Y_w_�GMu
�$�+u�߽RU�B�S	E��؍6T-}��.�U ����	���#���O~�ĕ�\��� ���וϤ��X�9����,]��G��Z�#�^�W��Y��g�Y�J�a���);jF.���tl2*�ڗ8��-�p�c\G:i"!M����RDI��Q�2�?g���	9jv._�UR�xd�9�RA}Ne�:���������������Y�9ՙ	E�5�e�i2��'�\���T,�6���9�r=�s�X��hG,�:;��hŊC}K��h�OE2���F��.[���H;���#�����%���n��/<��z/���n��Z)UB�4[4��w�<y�\0�l�R)/���z�O����ٳ�~�M�3̚y.���@,EI�c�Ci���s�{�l?��E/�J�b�d]O�X���s�A� ᠉&|[-�@ZQ�t��[ ]q���3����h?�/�_DU]�>%Jn*�5��!u�t�N���0���c��t�\��%�1���`M_�P����E8�BE���T�T��(,�!U+�@�R�L[�̯�*��&����������Ϗ^5��G�\�nnH%Zɮ���F6�6r���4&���2�_(Բx*K�.Ja�ݣ�!�oB&m-�
&���z�M)
Ŕo�p�e#��h@����~Q-L񘏢L5�����%H6�C	�O��a����Ae���F�1��Ѓbc�I�4(�]��J(|-~]m�5U6I$j*\�{��
�]��\1���}�V�5T�@��E�WL\�f(�O�'T$����DAM~/������d��
�B���%����X�'��C	��h�Bѷ3U�#�{�+������Xkʚk����^���2�&�,APUkCǧ�&�	9&��+C�!��z�������D�)R�f������@\Ǥ�]v�}(����}�w9"�bF�j�#Q��DO�\2��V�E�{&-�+ҁ�5xu��.�DR+���%5U5ITd��`����#C�E��n{\a��|��ƲK�c"�� @=�
	1��I�Π�e
�A��EKzP��t��&�c&�{-8�g�T�/��D�!�5[�*��\-��k@��HR��$��Mp�%<uYkM���Ր.��M�Ö�,��8=��&I3@^X#fH٦��{�⊥!��X(H��.Z��U� ����wLܔ��&���r�o�x��f���<�P�O���߭���7�^ׯ�bY��>�ip��&�ÇJ��W_�އ�j�qݵ7����/���7���e�Y�/7�KX6���A�\���݅�؄�~����b�Ҋ�*�	�"!7� X֯]��HȦ��P5#L���z�o�-|�t)F$�[@7��dow��O;�����6�Z䜃��_�<�W�caӭw#c(j��Z�;�Z�*��kxJQM��Q3Jv �ӷ�Ɗ�����n�G��w/���p�_>_�9��%6�1��? �~)�T���8�U�"�	b��S�ֺ�����9ˆ*Jb2�*��eC����
�`UԱ�ȇk$�*E63�o0M6�SU�����I&��cujf�S��9I5���U��j5�j&,:+�r�K��6�n�T��8>pK6�Zp� &�V�ւ^m���a��]>�$0~@�;RUKb#�Q�ae~*� �W[�JL��J�P��TU���"�g�%6�ߋN��j�"W�|�o���x��6u?��c\�C��\U�C�:��j�* ���bM�_#�B�Y�C!��@J�k�a�`�g�����6U�a(��k���	��sܨ�,c`�
����$ؓX����*.T,J#�5����MDC�jS��Z�u�ڤsTU�S]?���o8&Iʚuk�,\02����%��%r"�#�v�Q�&���9B[��E��\�������G�,:O�0�h�J�҃�XL�8��5KX��H�F�q��X����d�T�!떊��d*�	���o
%�	�X�f�#��Z2-�RI�D�A΃��������u\�F�!�v��3$)%#8�D*���T�"QT�Zr �M�TCJ�3��o����L4YO�`�p]=ݢ��w]��v�#g|ΏW����K@���q�7K����O�̇F����dǎ7��n����������cٺ=�(��GϺ..��j�1�}?�Bf�b6CH�L�˦�Gp�G�œ�B��`Rf�.�d��<�u=�/(�h8��(�!��X�"M���h3~�m�F�]��P,�.x���c���^�ဩ�s���cv�Ǯ�8b���V���sH���e��tg+�R��/U1c��Z Gfab�*��&ՙd�����D+;P-22��l����~��ӏn��\�W�~pꜯ�>�&Ot}V��.���[
�+�&#���ϕ�#j.#���s"�
�>M2q� eӐMI d* �l��4���B� �����-�O0�M���3���i~��b����p4F���������-�zW2سViH��M��v
��M���� uJ%��X<�m�]��@*	�l�� \�C���[�u�  k����ujm�Z��֢����ֵ�ג�S�ML����$Pʱ��,�����MX6XIT��yW�[ �7���W��d�v���Ājmdy�$�0Ib!�\?Q�y���Z�>ͦL�S�j����&ϗ�,���\�:�8�.PX���WQc�t.O4��u�(�(k�{���p4��t5t�.H��kǣ.j�9g�ze.`=�YF��/Q)��S���BјJ�="�uͯ]�&�4�S���F|���>���A<l�J8VEy$��5�s�¤�b���b2�ʰ�&#�����?��uv�moVu��/Tp��ڳ$��	���Q��.�̲��#�/��9Q�IK"�Yc��J&�%| �rs3̡6zH�"H�O:DrN���\�*��� H'��e��{��E��/J����PDD'������b+� "�����k��h?��׬S*��R��&{�ٳ����U?�����ܲp�巼��5��(܊I���ڃ�z�|��S��i`��r�<��#�[�-̜�&M`բ��t�-dK+H�T�*��@��6e�JGC��ϙ���K}�/Q�Vu��1�����.*1�(��������ڴ�%:�T���K�d
,L�W,��.�kk���^v��>z��}�yh-�)��tD�kn�?S����.U-���Z��QA\WA\�55�A<՞��巈�\�M���T!�|8��v�?��/��Ƴ�X�w��|8���H0�@[2Jf�<J�kGU��|v&���2����JU���b�i*���Z��*t�E�a%&�f�u	��7ⴒKmTՔ
j�CY/
�F��(�w ��;8�4�q���c�s-�ڰ<�~$%=��h�ɰ�z�>��U���m��$`��t��r�P�I ��j��Z�%���R�8	�@+�kAAq��s%!��#�����|�jŖ�]ZܮMD4���U�J��[�be�\Kj(�Z� ���&�*�VY�٪2+���(����d�1#���<�f/��R�Q����,�XTϯU��j몁�R��W&�;Y�����A蛆�fH�[�Y2���(J�Q�t�"e�a�ﶿbM��� $��Y���>y�	�)[������ 3gMW�#7�9�U��j��0��bDL�j)y���>l4
V�D*J]2����) �̓M�Hup5u� �=4���.;�&�A�wK��*�
kF����0C�ˠ��8�b�

5r�	!�ٮ�ֶ��.�|�Υ`x�>`�?j"�Jea	fB�p�d2�����B>�D��s�*��c�pʂY��@@��|gU��iH5�[q�V@�{#�v����ܩ���O�\�K@��3s÷˯��o�\^�oH>���U��c���͗]��s.S�3�̟~�I�/�O9?�}�o���rѬX��/�F� NM�*ʑ�s�^;q�6��/P��"��Gjnm��R�t�.T+T�"Q!�,F�ۜ��y��9Z�y�o	��F#��sl]�o�v���^���i�1�w��K�`e��#ܫ��A2q��d�o���k����fU
m=��s�2�
�JAo��}����?�;���C��;���x��G�����FkrA�C����@�-�X�+�Y��P@m2MuuJ)K\�d�L[y ˊ����%U
th�U��VY�nes��,��W ��bx�߾�*H6i�K[_�*պ�V*�0l�`{��Ȅ�c;�U��Ͽ�D{{Mdi_��B�V5��P��be����-o	�R�*I��6����e����p���R��k�fm�4���g�*5�%q_U�vu����/���|�@8R(z����K@w�
����1�Z�FmЂ��}�j��uu)5F
ME;��y9'����R����@M3��6IP��b��R�y~ ��@}֡$�6���S�d��9�$S� �bfP%L��Q厍]up=G}~Il��J��cL���@T���IB#�]���Q�=J�"�HLU��g��];gr]���d�
��nI0j�^*^��X�ٳ��
�'S��%��.�1C�C1�#���R������1Z�a^{�eF�و�c7e�`���7_�"��X�J�BΓ	خJ�%��Ap#j�_��x�{#�mx96r�1T���ܗ�m�(Y%R)߿]��l��>����}j(��F'r�%�ƅ�ԘDF�*��Ð�揁��.�OɒL�l�����]S3n�Ĭ�l�y��3�8����O��K@���u�K�����^��� _4�PaD�������$@��P�ڇ����`���Y�ٗ��)�M���Ա!UۣZ�b�eZ��W��Qk����9�I�y��pS��IN�б$i���xn��VĬO1j��<������[��>��M
5�C3B���i���g�����æ2��3�1'e0�Q;�d��R����DS�
,&�B� ]n`���FS�u��I��L�` A.#8��Gs�%�PM�,��ֻ{l�彛��!'���g�䢕]���ݻ�P    IDAT����/�;��)�����$�0A	{6�b�X8�S���[�֟T�R���'�(��Td��+
{RQ�(0"�*3V��Y�7dL#�xi3��V�Q���
�RJ��[ۮJ
�|��Tp�E԰�c�Mh	�y���a���ω��3Cɋ(drPװ=����F͓�+�T����b�xOU�~���#���_��6��~9����d�S���yPsXWh=�(B�ۡٻ*�U�(-ti��	Gm�.�̌��,�l]%��� �x�2C��Y�SuRJ�
����6��(�!����ķ[��rY�Mm�Bw+U0�7��G/�V0T3SiY���*1jM�P�I�Y(��Tw"U,%��9\��:���7S�,Y�����Q����] ��`*���B��*p���G�����������K��$�:k��HO�]_�^�=E���X0��7K��9z�`<Nɵ�TK���!�s��1S#`��kۉ�,��W�z�P��cN=��+��)z��B�
V��)|��4(T�����@�2�j����|i�P�¯�kI�\#�4t���Mf��8��������1
�R��p��&�ʿ�k6{\O�4�[H�V�A]��hE��7�jG#6��>�d:�f�Q�O�~�V�!���_���8�W����>�zV�لm&!g�@��u�J���L��*Z2S�d�s�n��jl!k����12��j9��8�I=,Yx2���e�1�L�kG�}�_��o':�B�G�GT��%���i��1o~���F�屺o �*�V�A!5D3����׿ޟÏ<�cN�A�eCʂ��l���ف�̃Q���/U�'��AH	hU�'dh[eن)���a��u�2A�B$��=��uR�\ƨ�����QYֹ���r����T㈸׶]��R���WC#y�Ћ⦴�="r<z�r4FlU�Kr��.H6_Pv2��u͡K*�T\Ǫj�[�NIK=�%ɏ)�[o3��6ڈ�^���Rh�TQ�lW�$P����~p�`?8�%�`e��n�)�,���U��b�=���*��H�5���+��|��v��2�ZWxh����qKE�*���!%"hc��q|D�j�����z�C�`����Sc���@d��x�E�dO��\�$�*��H��Т_.�µV�<O���5����/s�r���BA�
 �>�6��U�
�^u����P�(��z� ��[M3u*U9V�H�)����P#��I���\�2cU�_u �j-�$�U_���H㷿�2�@Z�~����x.Z�P�1�[�r�8�n(�\z��t���� �\�H4�A�2Zpe��b�_��@Ύ��r������w��פi��A>� ��$'����H5�{�^��#��X��/?S��mvݛ��F�0�"uXr�-�$�*W�jɆi�a�"�q_t<�GQ�[ #Yw����J��D�OX�����oJr�IwP|�?)�X>sA�5*�����ߑ�Q��M�t~�$XX����c2�J]�Q�Hz�ؚ���%$X)��؆�^�6����c��u���O��W~�{�}����lPV?R�r����(���k#-ni{�)fz	U4xi^���;u*���n����T�+}OlAgF�[-��F#�bL1��)4"i+rT�e��d�j`��]���=��`����{=U����M�(045�}���o8y�y�����B	[��֢�g)�z�!nDa0vn1G2Џ�
��ށ~􈏪��U�K4+>{��Ta�@��G[�f������wӧR�&��~��|���X�T�&��i�c�G
	S�<r�]�#.���w��)�pW��џ-+@�l֒\)Nx�����uS����eF�h߀R�#�<�\)˻�z�P���)����`�ۭ��~{���8���eG3]�n��nИ�iL��\�X�iZGl� ٜ�|JK�&��Rr�d�2��L� f4I5_����K�6�P�|0�\i����z��EUG�+�:���#Q)�H;ZpvEu�_1N3��f�9!		�&]��P�%Q�j��@���N$�@�X�0K��|�TI��9�!Y��� �D�(1z�0�~�%�TTU��#@��BGK>"��b�H2S���P��l�ka��⊚V��� �,�JA����t�����mO�Pr߱�*.LP�L_�A��l����xU�d�nTl��eQ�N�h�A"�T	��>OC��R�b�յWu�y�Y�LU);Bj�d$�5)S�:��` G��y�P�jI�l�W�C�{�T�s�Dx4[ub���J�BpC[:l��U+�j(
���E�_^!���UJx%�8��\�r%Ȁ80�6Q���T{��:v�/��4t|�R��8��r6�4�@�𩋧��.��*_wd�d�ʹ��$t�x$N�����h>��p�}�tɉ N�T�u�H"�q<�L�"1a|��#f���0E�V#�ա�|�ga$äM��Ѭ*;vD��s��G�����K�R��ġ���u�?�޷ggq��	Y.z.���N�X���I���'��M"l���aD��?����΢�k0�!�aAq��bI��9��q4���c�4�u:bq�l����WҀ�&��QVw��>;��cm֡+[ W�*t� g3�*7������*��I[l���ſ�M<�!yA�-*傯�$V����f��[�鴢	�n;%���ٯ)�Wb�U�R��B�T]�u��|������9jjT�Wq􁻳��7i�y���3���8v�Q������П�7�$��l��,��X�NQ����&�?|��O��C����.��<��3<��+T�0���Ŷ;���`)>�C{s=�R�e?|���Mkc}��ra�p�T��f��vg���{�m�a�m���ǹ�ɿh�h<��	���[��,R�6Uzן�kA��
�k��#�!���ƠC&�$m�4���V�� �kl��e�R��(l��*��FɊ�iD�;E,C�&��W	��*`U4V���.��z���tP���a�l���������:'RT><����1�+�ۜ���8�F�%�l��t�.IU�K�ʦt!$FB�'ObѪ�t	gX���"�)@��4T�&U�c7�R	SE]C�
bNU�Xb8��6���T�>eV��j��x,�2~u��T���!�AV��a��+ʀ` 4���pu�I�P�ձ4��|�ҕ-bF#T��I���g�����*Q*����"G�@�NY��Iԫ��IR&#�X,ze���~�:����@���$�r��4�����0�|�H�ZEGuq�j�x,L_�:o����9H_M��%��fD��"�+3��h0hy��%(�����{<�Pt	'�X֮�ahU�F��:VY���0�|�9
��$Y,R�K ��J���b�-��K��Z�]B�8U�fU��>�(�فuDR	�f�*a�Hf,N�RP�Ʋ|�G�.H�p�I,��:��}��v<�,���藀�w�{������0bJx!"�ځ.���|/	�,|U�K2k�(�s��p��~��w^�����5�%ä����9Je��(�*Jۦ�.����\b�Kz}'T*���ol ���;�
cD��Z�IU2�`��\?��]Ru��ժd*��e+Vq�3v�f�{!#�L�T��*K*i�e��2+Pc���d#U=�a��J}�v�6x�N%�"ŅT��e�,��������Pe��6��/���W��S�q�q���[��O⏷��_��H]n��P��=�;��^y����l��$�W-��s%'y 7��r.<o�_�{�x�n��N�6�՟a��Id�%/Z�6�����]d������v�T��^e)��v�C��j6zٮ�_Ǫ>�h�H�TD���%�H�u�he<\��$C�Z8A�,O�T����E�r�h|4���j��+�����n!Ͽ�Ol�	=�BZ��ef��L(
���.
�F@h8e�!Au;dm�h��*�&a4T���1��׷Z漭��kM��5���\OW�D �D�M�hC��h��fj�D�����4m�M,[�I}k�
����%� �r7��ƣ���"�sy%��xMv��L�֨�W�R�K�[*�y9EذU'�w G&_%o!�'+A-�Dd{+C:8E�luQ_>W���:��EaB���`���T�K���$U+�.�FWZ�B��G"�dʿB��xϮ2��@(N��v��y?J�J�oUs*!�h�Jz4$�v�P�����V���wg��� f�Qͽ�}L�r���x���f�I��%f�U-,-H!���
��8(p��<Ւ߭1m�E��e�=va]W?�#I*Yhѕ,�`_���m���R�=W�U֒���S�s�+:��dˮ�L�b&�|���������.�S��*�66�R���kh W�1�-a���8�Eaˈ��+;W��˸��]��$�:��Q�vv��@ RG�"vYSM\���`��7������"+;s�]�Út�����U��%��^���Ib�^���SG�os��t�0�����/�'��o}u׋_/��	ב˕�T*�Pf����;�`��ő
��c�r�D4ΤM����.��3��[��M�L.�z)�W3��)���j�I�0�D����+��@%�
��,<��2�"=鴢$	�C�g�*��i������60TKx���<��#�u~�1�v�Ts_�rq*2����5|�Jk]T�sݖ(8QR�&���y��+7*��Q�2�t]�~s���޹r��1�Y�簺3C�Xe�ؑl�I��s���6�Od�_o������O?ϧ_|�e{jƜΖ���ִkc��.J�=kW�jj����~����Iǟ��e+y��jhQ�~��Z�^tSC�]�.�ɥ�8��l���|�)�q���X���n2�֭P��w$k��o֪�]I0g�ADQX�cOݭ<�g_t#g^x)V����#�BY�(�����D�'�Ak�F��������~�UYL���Ό�o`Yw�@[+E�W��͏�~F�ֳ��{�f�j�y�e�u$眶7��d���{Y�.KIo��D#�r^&�8�~�����;mK�`��?���~X�6ї���\�bڌYD�G�a���"�@���jí�������=lwf�q �^�(_-\J �δTG�v7gL݇��ی����]���{<��X�z��&�}��w,�*D��f��{��v���8��M>W�9�Ҝ���۸�8z(!1]�Rn�@u�I�"�8a�
�����N�3��(Xp������`��k�����.�	�2c�GL�E���Z��V���l2>�Ï��󾢳{��-.u�RE�^�d�kz
W�檌���g�ӏ?��|�1G©�Ds
��������e��u�d��:��˩G�Ǝ;�̩�A&��н&3k��4Fa·K���g�-k�C�5_!k���`W�l��x��`�#p����u�V����G^bm_��:�p(HԳ(��d�7c�=�`��Kx酗��װ�n,]c3����$�8��� �6�Jصp����l��-�(�k���.�Wn�{�����N��x<ʰ�!��(j��)�KP����p�T�:eN��A���'R�N�-N��� ��.~ҁ�p�h�H�JMq����,���^�r1FC+^�$��(li�RlQ��Vaǎ��sN�q�����|�_�O�YoͿ�Ͼ?��h#_�	�sl��Cw�X�ן�C��X�t%]��hood�����hI%9��_s��3�aMAe���pi�'�Y�n~���.�Tښ�ɉ͡�D��[����"!�qHK����)�gH,e	�pCꊡn�k�����{�QrV�����y�wl@:�#�3j�xF������u\�����������9�ݕ������y����Z���U�9����e��8t�٤6`�7������7�ﶛi�kDwJL�tU�DW��{k��Lmꮆ���Tfƛm�9_~9W�;��9��Z���P֦L�D$磏>!M��]d)͈���b�ɬZ��r1����<@ٟ.]��c�;^?��cB����dGO��c��ڛ�;�jh"�����~�7���#|��;�p�y�gY��f���n��&)�!Ҷ�v
�����2e��<~�q\|ɟx���T�3Q�W��?�'_�R��ǥ�*�i�K<q�L������|��d��2|D3K��L;���{#�J��2@<��)��&���G�P 9�V�����#�ǧ�|�����g�u�W�?b\bJ�e�+���jq2��^���n��3������>��:�FJ%wpS�˟.;F`���\>�r�jun�����d.��U�z���j�`�3�\���ҳ�s�A�X����f5���`���(Ͻ�=W��0n�h���9�A݅�
^��2�������~Ťɛ�+��)����soeY_�P}���V.�4E���*��"FD�e�^	�{9��9��&%`� ����������|b�F*z'�LƲ	F�XT�z8���̭��[�Y���O�V����V��f���Qg_�@5��A]@��
���sו�s�A۲�N�1q���x�=�l��Fq��r�ϩ1�-�`#�.6����7�MG���z�i�Z�X*�͏|��D�iM�]��nv�<��g��:S�d� �����W�ٖ#��xO��`�D\w��]��zf��N�]%nV7�p�%��Gsx�g��ܥ\r�]$G�}��A+�h
V�x܆T����W$蕨�9��{��8��[���CO�䉃��i{��_l�{f�D
X���?����=
�p���em��ut�c���5B1Y�0��FRxV�m�ÿT���$�g��W������|vA!1\�G��>v�s��v�MC��V�D���_@[k�rY2��Zѝӎ?�U}����ɬr��pݫ�ٶR��o&����D����:��S�",W,�!����*r�ȗ)Do��ShT1���*���O3s�9}���)ۃ�,#��H����o9jCƌ��[� �k�|�ӯ�~��<�b�2�;�0�ڤ��������2j�(�V�/?�Ƨ7���1O��!��t�gy��3�Ƌ����`d�*�]��E>_���MoQ�2��jIn6e���6��r���\�b�J`�� �Tb�<5��U�lm�P�R�#gժUy�<��ÄC��"�<^��[D�>j$�]��
E�a�vB�u.��z.��>�]��hc�R�
i=�x�[yw�k<t��t�m�_��}���aC���3y"���Z���Kg�v��zԎ�ö��&�����y����q�z�Ϻ���q�=�Gq�*�j2�r<W]� f����N��1�s��aGr��'rЉW��'L�e$9���utw3󴣹�艜7�b�Z������)-�|��u��ĚG��	��5o�����7�*�����ho�RYf� x~���<��8�z-:��uXn Sj��r�|�[C�Y���7݌o�b�ܹ����r�m���Fr��b��Ò��k��m��]��؍��v	W^4��aI��Yf��N�M��!���g�ƻ+�ئ$o�ji��<�ڣ������W���ϟ��>�pF�ِ��{�c/��y+�⭊-��P@���oe�/����~�8�"��(�X����E}D�Ow��Ï=�m5��|�i'/��*_|��\`F�I�#�5�������S��{�擹<���\p�<��\v�L��r"g��E>Z�
]�V�����.ᶋ��wf̔�8��c���C���kY��w\{�]��9��	��:^����p�U���[X���W��g2ݜu�����������nV�j��fՆ�U*��9��9�ĝ���L��5���������9��~s�M���G�w� ������kǈ�F���vb�&��p$�o��m7�ω'O�O�s���5���D�%~52�7���lV�H�(���jX紋g��r��ل6վ�
�����-y��L�)�d�ܯ�����k���v�]�m�����j��}:�t�Y�    IDATG�I)�������֩;��
<��b~����]�������HG��D�g�a�9y7F%�dY#!�MVd]KRY��>-�R�p�ʡ���J��|O��t֯&$s.�JjQ�w����*�����T�pK���$ ��f`F��҄լ\h7%� TE�����j�jΜ�;f�<�t����ս��5jC>��F�è��J\C@P7�����&���H��g�*.:�7d���wߠXʱ���������3b�0��^D$Y���$G)����8�]}��M�fݥ�-AO�z�U]�L⥝�E�Xd׬\�{�����*������0�|���+��´��(�O>��H8��c���7���u���|�ŧ���R���t�%[)��v��?�E�$�r�-)�����[���X��#]6��s^���y�ٻ?z8�~��ͷ،�3Ț�>�w����o�%;�D�<Q�B(lпj9�s ����uucF��[��SO;��?X7ߏ�2���<Z��]Ǐ����dֹ������ܗx��/���YL=�μ�dθ�.�Y���7ba�ф��q�IGr��M�v��qC-��s���q��;�eX�.Ǟ��$<b2�)NdN.Ǩ� /=x��<+W����D�vӘ�2a�8����jE�D3%�&�G�2�\��l��Hf�9�|�̾��S�P��c�m��k-~s���b��Y���Q��G�cͼ%\2�,�L�_���[o~���ϼz/7?�,w��5�a�(�Y��0�0"T�g/��oQ ��3�P�C?�޾���9��_��@�C����4AS�� -Q���#hw�UiU�^	k�
���vښ��~4�`�c8����y�:E�����y���p��T+y� ���[�+_EG���˩�����^�g_�k�`��[p����G ~>�Q��\�m3��w���e��M���)'�Lתu<��_1�8�+�	Rm#�fi���%�8��}8���X����Vν`&?���K�&5r2#�m��ZEY0��Ws�IGp�;p���ITx��������w�ȟ���[n�oN���jL��=��U���i��p*[Oބ:]��c�{��v7"ax��e\y�C8�(���!RL�u����\��������X
��#X�b�1��p�DN��n>XY�N�S�\�Bw��0�1��{��g}H��A�;����ƣ��*QE���+��`<F����ɒ���ZF��4�>��ض#�ޜ�v��ߌ�?�����t���]������?Ԅeċv�#�axR������Uf����3F�v����e��Y,_WPS��T�XZU����L��	�ZPQK��$ҥb[I���6�;{}�϶�z�{�/�Qq\�V%kWK��v��j
0Ӑ�c�5�t\s�"oN��I>�G�PT��>��1c�Ғj�S"n�.���H�F����1��}9����^A,b��?ͨQ���U�ʰ����{�?�|43�aF����� A@���k����)|���4�ձz�J�<�Pרֱn�%_�P�������>g��vTh����L�2E�/]�:�uqE����r�q�х��7�d�/RZ��Q�G��i����������t�h�b,-�!G��9��K8���Y��kހu}]����Z~�����h�/n��R͍��zn��qV�$|Dqɥ{""���\�o�ۉ�O;��S�r@�F�bH�6��}�%HuP�v�Q ��	d�y��;�T<N:m:q(k;���'�����㙰�A�`F�S1��d���� ;M�����/�5�>Dcs��+���i�y®|���*����IW2�'[�:�l��]��������TB(V~���ĬY�q���XܕCFq��fR�_�~[�f��'����~��իhL��w���6��7?����G�q4%LB23uD�t3�=�Y�v�Y�l
p��౧.�ϯ|�Uw�!�1��Ջn��з��gNe�>�����s�*#�ɛt�uY���+��=�T���H@��,%�#�N]��ٺ���
a��ս��<�'ƍ��PX�J�����)�O�sOf�q��u�B��� QI���]�r������rR J
<��w\t���*�rI�ʾл����>;o��y��~iW\y�J^_x�:^~{������,����%B��Y)P��fxC���>��'7���[�yW�O�c�b�#&F��F��c��$�vs?_��w<��;��w�����fM���G_H�m#pe�'�q�}+9��_1�C�}�;�1�4��]���gO��C�慷�̺�f"��?�G7��*Y&7x<v�e�x�k<��gI���P�_��sfpԱ���+�����+�ri���-��%JBQ4B��z������g�{���S�1e�mx���1f$F}#]n���$���<�3?y{�������*��W~nk�Y���~{�_?Yx��jW�B�^���'�B�Y�j�J�@P�*6�>�+�R-�r�>�ѓ�(��!z�)lpzӂ-�lLQ��	J�Z7����^��l���5C�e�b�`�l��x�M�g_�zt�W��Q���n����z�t~�ժ2��=��F'��;�����&��B�'����G>�n��6Vt�\�R>|�Q�b'�|�I�N�<�_��Fҽ��ށn.^ʷ߯fMg?}^}�%��ڋ���ˊ�\,hmoU�A�K��p��B۪�������V[m���z��T2#�b�)~��H���S*+<�}�N�V[m��E�kK�4v�%�Ɋ޶����ׯ���W��v�}Wu	�=�JN>�z.�%9�C��J� �]V�� ��&t�`���8�tR�ñ͸�߈y��H�.�,�Rʬ%�G���N�P0��4�*�#�8����-cK��~��vs*�~����[u�4���=��p�]���>�ͬ��7�������f��|21�H�����Y�5����s��nN�*"5&��:��$�u�d�w�0��5l��a������=��ނBL� ��YG�03�8|�9h���.��v���/�篯S	7㆛�� �%�^�l�1��=��&l�E���O?�1c�o�ԩ;����eP׫�Ţ� �`/�cEN9�P]�{凉��s�9KI�>��y��Uh�f<#�@d	ښ���r§��o%%�A��+��A.��5>��kH5��2GW㱪�,l�b�1h4����Lޠ��/��(�������{�/T�mT��JڅKV���K�S�N�М�?��J�5r��G��[�d�nH�S��0#���$G��y�B'�s��;|���z'�@)`�)!3��ԙ�t[Lٔ��N2������J�p8��z�������0,�P'n��L��Qf��擹_+��r�2z9�yg����"?�"�p
�Q\�DL�R���l�d��˰�g@��h�
�@?��c'��e{n��~V�L�h#��D��*�!�`E�a�B����y��|��r/<x/��7=��r�]a¯��='1�����#D]����>y���	�?���Z̃?t��Ϊ����J���<<ɭ���ؘ��:����}7��F��҅�Y�vg�u2�^z)�� �hduO�r���g�_m�╫M�ڄ�d�-�sщ�/ARG��r�<��a��7�*�X�%��4�����5K�9�L:K�RV�2o��Y�e�^I{�h�?�|6ؠ�1����8N�o��z�w$��n��[�^'^A�y<Z�LGc�����q5�>���2��%<� �*�T�-(Ӷ�-T�b���>|����՗TU��K���J%K��d\ <bq�����6�̙�>���ڵk��*0�U��|7.%7j)��	�ƫ��5�����.]�:�=b��vS�y���'��J �;�f�}�U:��9��vK���0z8��4�fS��崓NaՊ�̝;�w���[��p����?�`M_��!�cy�P���d��x8��5Vf=!��t,��p�_��K$�=��5������Y+K4���p,���3е�hз,���&,#DZ�J�P<�;؃[����a�:1B8���U*H��6E#��x[��VY�ߧx�f�^�ȱmH��u�𕻂Mh���D�FT_��������4]Fv4�nm�L�E�:1��cĚ�t�@T�f��{�SN���ђ���4]݃�7�����T\=4=��J¹wM���b3�	�Ȇ�����n�o��${�BDD�\��M��hU��r�})^WxM�`%�$Db�(�	q<,P3/H�*m����	7;�U���1�
K�oMz�b�۰�W�>F[�a�#�j�#>馺���0P��[�.��Xa�'�k�7���C�hlk'k��F�)�Fi
��Ŕ��c�_��>���:�m��%��
*�*��C$$]�8hl��_�w�Tu�5�o�P9t��DD0�9���1+��QA1c�1gQ�4**�9�� �c�T]�n�M��<���}뛵f����a/Y�Mwu��;��:�6������B�௢V`oױa�<��A�2�ydSCO ]�t.��hޡ!�?7X%��pL�<v�̡�-�ԣ�:���jq��
��y@NH��7!�'��q��o�q��U(d6���8���T������{�:�{��P7�/��9-����Ԫ��e2ص_䳷��4����_���!��t���#�|��KmN =�y\;���3�B�m�e�J9,_�
�}�)��2��鋝�M�ܗ���>����������	�YO\��L6�`4����A��̦��j���zGwj�b����,qMG��w���c���uD#	,�f�F�j��&!D���G`�ڕhjnB�������I\~���<i{�=�53�	}��0�N��ѣ�`�}w¢e��	����T2������V,@Р��!����	�2�|�F���:���ƛ���O�����:-Uyp��m�SN��b�X���اY�3g��_��W�p����?�����Џ���dhS·�ۋ�o��U�2e
>������"���0sEIbb�]º�;Q,q�a� ����.�G��,����Aw6��d��V���wx��g���᥹�����g_|�~|��{+>^��Ɓ�s�o?�b�(��N��N�j����h�ĝ&��?MD���଻�Ŝ�?B����W����GJ���u���ɹ7��yDC2��´�~¯9��P�c&��EDA)$�/��e�aŐq���e\pʋ�
<�,�`���(]�Hh�b��6���#�E��RZ�&�@��(&^�DCU=�6���>����/�����m�A�h���f�cƕ��'^�XO5�@$V�|��Rz�Q"f@󇥀�6#p5�܊}h�|�rJ:5]�fٕ�/Fx�Q��/�e"�4��l��=��!?�f'��4'�a������ǌ@Tȩ�S���b.C���\�mT�ն�5	���o�W$Zy��+,��@���V4?4O-<�+_1��;�l/�>���(!�L:#�%4)\��GN�$�#��a���n�n�k��b�Q�N*;}��a��9QԈ3<��"v�uG46$��S� ���G�U�'@v)+��d�?*�Hq���cҲ�JoyehA*	�"�����MJjJ�qljY���>}�����1p�x��i��L��
�JH-c�Z��&�gV.��k�+�ú�x�'Q�M b�����O^{W@�����V�S��Q#T3�I�B�}�N��_���K������؛�Ysăo�R.� �5`�r������nї����P[[�|� ,Y=�`�j�Qt�nc^���8�1S��&1aX_�ߞX�b	��jźtя�c��s��6���!O&�H�\TG����ǒ�2eNQ��K����T��N;MBs�Ẓ.ڈ#���S0l�p�r���H�kS��F�$:��tR��	s�h��mY4bRe�}�M�*��Fr�D,��|��Kh���$���3��G�4��:9^En7������G��G$Bu-}�K��"��dSG�̚���������k�a�̙x���Ň��5Q��yQ��m)�Dbb�Ai�䉻�d������/��e���Ć��PSU�D4��-F<:���!��n9y��G���g#_vіLÈ� ��/�	�|��y�1���G�;�\sí�����O��o��:QT9AJT�hW��m��z���DsD�Eg�������,�=�<��%��fd����yP�by�2kݣ����t�F��W\y)�۹g�z��@�U��a�L�!m��<w���/(p�m������8�[Q5�U�po��:rm�Q�6u�*B���g�|��8�ɸ��y�~I���(B�ʰ2Y�Ե�My��rI4�U\sͥX�كf߃D� ��X���箉���[D�i�C�]��d��Fx�!(�i�"dY�,�>$�Å�^��v�b����Igc^<�e(��U��X�hPc�l'��m�#�C�_zɓǩ<������E�W�J���]Mr��m�	�|l�� �`Ѱ�� ��7�������m���w�ކ�/�1�������y��8���7��K�������3w��'?�����'=��)��@���Ɓ��"��9�4>t��çy(XD�ty����<�.G���x��M�}�v�y����W�����8|�+`�H�ajk�^�+�6�NII��B#Y�2��4R�_qd�
����@1�0����G�綸n�����[-����TUC	G��Ӄ��Oи�x��&A��(�^����X���濠XA�P$ɮ:��X�b	-�M���䃥�z���5�.�������������5�<�޷��Ț*�t�C�;U3D��3����;��?����D�B6��ǎC>�A&ۍt����:��]�c�õ7ߏH8�?�3�������O�D2Ջc�>[��o��O��&f\u�$��M���?�"�;��y�lhA��t*��n�t��/��L08&�H����tz���鸔�f�D�"��$:�$� 7��ɷV��ۆ]&�Dw�O����TB��I�F$�k���ͩ9���y��>�f|��<|��'B��i;�Vo�� ŗ�,�]=�o��Ç�W��+���/�SҘ��yˌ�,��aۚL�N����nL�u�H�8��2i"�~�yī�嗈NJ�tC'H�c\c��F�u�n=
��	qā�q��x�ݏ��۟!�8#Go���k0������W���_��ٷ��'�৥+��/��ヅP�w,&Nq��)?, Ă�m�SHڙ�Bo��x>�j!��}��y̡f�lEG)߃�9K94�C��v�B�H���B����	8k�CX�� FUVA4��i�*&TJ��DD�p�*B�c�������+��#),T>���B�������-�@>+�}��cO9g_�2>�y�xc�ۡ�r������.�%���CBup�-7c�ʍ��{`EF��a-�DYc��H��E��-��'�}�G�v1���p�j�c-�҈�h����*x�h���U��{�T����&�
�#q�f�w#�U��5�q�I'�Qbd}���YAy���D/fN���XtE�NB�Ϭ��n�����Cg����������/��	�����#�* �,V5�ir����PҭرI�\�s�z	_.� �f`e-�Y��P6P��wt�O=y|]�+I��N3���ۡF�J�D>~����AcX�3�����|���}-�$( �%�ŧ�#N��"�@���(�I��$�,��f(����rr|1���V��=���8i@Ktތ�x��x�/�D�QS����U��,|�4�-=x�՛����knE�ր�ЀVD�.���J@�
ubo��icJs��wN�e�����Oޙ�'���]�������,�E���C/��Hi� �մ}ex {�|Y�фF9���Iv"���]�ݷ��.<_��?�yU����tw�%B8����e�R�{�-�~�F�:w>.��z���<n#��cEp����ne+��|E��    IDATz�N;��p���J�� ����	�KjZ.K�]x����Q��d�z�G�y�)���Xt�ѱa��:�.����Gs#}�K��efOs�3��%���=w�ƼW������Ej�j�:��W�|܉��3��LJ�tN�ۼ7���7݄'�x���E����R[�(?�'�A��WEL�uW�X�Jnk�}������_.�ƨ�\��� _̡�����`����;��s
���s<�ĳXْD����]@g{^|�.l��t�s�r�����?_��]у��s�(f!4OaxMz�j{Ծ��)r�~��
���h�7������B��uB�R�"��87^~ ����O��y~�@��|���ՃQ�ǳ��L�JY\t�p��}ElQ�P�*!�e��,Y�Ɣ3��8Z���XJ*�1}�x��cA0z�GE�]8� ��	|��r�Zy͢��ӛp�'�=�m^�誈=B��0�58���3z�>�, ��lf�~=^7Յ�$�{e&^{��~���E�	BSx�B��1��<a��	΂��H�V�IѕtB��XSM���xJ:�X(����ɝϽ���ԫR�*Ŝ�;�?��Y�K��3ғ�#��Ixq��)l���!0Q�k����K��cN����1�뇉�sQ�L*�܍$C#,�	i�T+n=� �9�]yڊ:�xJ�{�z�	pqL	�-^�[���Z
B�
����I�&t��E%�'��͕���A��Y���p�a���G����vN��]F"�@�r%��S���"D�5�6c~58ҀV�R9 ����|����lfO7F7E���ǡ��m+�a�m�⫥K1uߝq�S�ṷ>C��! �7A�+���e,n9m��	wκ/=u/����?�0�&�>n��X�҅D8�"C�ؗU���=A[��2v�z��'��O����������c�+N������G2S���a�ڝ/2y@:a.C"u�$~�2m4^�
���Ɏ����Ga�b�}�n8︩�i]������c�Γp��{�K/G�~$>[�Hv���F�ώ�5�,L��$N?e6-[���|�P_,m�Eow>r?�nW\uL����BsVK��DQV�d��L�"���ta��3w�BU�
����E�:�m��n��X�ɫ�{��Cj�s����Lߪ^�����&jM�����'X�ӏp,�(���:t��_~^�!�U���^��8��������狉�n&\U���J��W�<�������{���?����}��gӕ�0Wݕ*V��*d,��D�c���(yY\7�j<p�CX�d���K��1��e�&�1\ۯ�����%��Ţ��ɩ��A��$�Uq�JW���$���	�ul�hd�zŲ�|*=P��.����@�$j�2̶8|��x��c��7�X߾��c{p����F�]p-Z�up���-d��Ȭ[���<�8��J��j����Щ���3�)'���6p�, ��1�Z�3w��d�&|�K+�@=���T�30t�|�X���f`��۪(lZ���O�����;��="�[ʣF/c׉[a�gkq�����3
9���Ⴤ��H���΢�/�w���;nys^�1�����l�˲%�"�3�O��(��.1�64ں2DI
�˕S�x������q�����ʴ�b��ÂM�"Nr�>��|�"��k�JR��*��؞O��P1�����5{pz�"�1�����C%"b�=M	"��vlT9=���GBQ�8s���D��ಈ���3�rCC��4o$��3�s��+ZD��d9*S�~�����1�n!\z�R���g`x���gc�S'T��a G;8# =���逪Aox&��A���d���L��B�W�	�ڭL"�G4̹��R�Eg����M�7�rμ�2�߱7>��}�D�Jj	�3Ӄ���iS�`�����b��ݔBO���v�|�W����Q�-%�B$�� �?5��KaJ���˞�Q����3����]��i��}�-�����I!g���-����y2))�^���U`�
l���-]k.�D\C�}9N=h2N>|<n��&\vɥX��Z���=��~�����_}���\A�6a�F\t�3����Qm _/���!x�ٹ�������
�x�9��GF-J�������a3�ȵ�7\I���%Q�t�xb�-*��5{���,��)�ߎذ�+,���jr�q�fN���M�-��4�?v�ר�Y3/��������%L�aG�4q'<�ȃ8�sd_�f=���� $a��f����p뭷��^@OO�t�g�~*>��Q
L�:=���j�P����G..qdUo�����3���w�=��%�f5t� �1.��#��#�R1e�=Ѷ�w��L��Z�
6zi�AoB�J��G9�B��
�R�@e��Go�tQY��QUC�L/ @�<،�պE�n�E#�x%�UX��B�i(r!J�22)��M�c�`�1�X<���x�7Qf��?�\2���_����3ι?�+B�j�u���9� ������a��e��
�+��ۂ_{
��a�coF9� K3e_kd<���ǎ�#s��·H Ȑ��8�}1��?��_Ʒ�{�Ǣ0˶dֻ鍸�#�Ϯ͘v�^BR$�C�����.��p���5C�薡����O�'�ew��+O^���w ��M������Fr�JR���3D�����/��ã=�}>I�@
5��,�D��aQ�^�l���2��	��TUijU"<z��e�e̫d��/V�����X���4��6b�	�qǕ�M���|�T������lTZ7��}.��Xh��Z���?��O����(:�L���86�n��WHg���ca�,���]�"��υ�@z���X!�r�G5���}�8�w͞8����8�0#��(��:y�������P�pp(� z�	���lq�t%�\�mѧ�F��D��uX���qˬ�հ��d�lX��Ç����/���Xۆ#k����sp֡Sp�a���\�(P�����W��Q�(5�f%Q>�����!��Li���);��O�����������������K��Q.���%0��a1��R�.vѳ�J&|�1F��p8������<��n�Ѐ�����n����:�,���5	�b�D=��.ַo�!���X�罉�>��z2��
�)�/���{���0o��!|�:��>�l�6��r�:T�W=�t��,m=�w�K�B�V��MDu���I�>`�����7���x(#���h@O�����)S�T�po��j|��;X�v�8�]z�t��p�5�����U3����?@(���4h �A��6���:<�У�nͦ�x������ԧ{��O�I��ԭ�nh���Hj%o�=���
�"�|�q����$g��c���$�6�B&ec�}G*]���ݎ#�=���H�5����E\��#���������oq��Y���pڹg`�-/�ïV �H��D��I0�ǡ���a�a8�W���.� 5�G������8�/
���y|�s;2�ʄ/}|e�[��k�ѕα�����v��#�A��E�>��Tz8^���7�Ơ�>��-X�lɑ5�2J�4�}�{�uˣH�Bi#T�EЦ�u	Æ7"��A{G! ��^L�4�\x���R���S$�-�1r@�$����]V!��̔�C���B��x#�}�)��MBh�$M�)L��ޚ�~���T�W7���G����߼��52�Z+�.�G����O�s���q�f������lN�dsW|ι�a|*?���}�By_�""M�<�sB�s��=������U���#W��@�~6*JYJ��q�`SG7:� ٸ���I���)�,q-���@d�1d0V���#�!u�;P}Y8Ţȿ,:�����*�Dmȇ|6	=B�ѵ�K����C�~E�� �ﻁ�?�T�F�_�L&���,9�$\hj .�9�-���x@���'S��2�ƄrF�7��}�8�<ρ����� ��pӅ'`�m�c��9X�֋R�����lވ��H���Qȷ.�e'��'[��Y�G�}�q z�h�姑�n!���IF9�=�x��m�����������'��w�������Bu0-�M☉�� ��,�~ѫze>ϕ���qrB�W��5U��X�\2�6���}�&YE�(a!D�p��$��)dv7�VK�Ѳ��@�dq���QP�x劬���aD�)���q� A��͸?�?!��
�bƲ#�Ra�����R( �Ҏ�j?�w<��v�'���"N�FА�v���p(&Mĥ�\�/>~K� �d��K.��mv��3g��+/��s_śo~�澃��ى�Gb��!x��9�5k{�q�������c�⵹/b�����v8���*:�~?��:p���⫯������/<�|��T,�;oÊe˥h�x�	8���v�j ��;NF�_��N:'�w5Vv�U7�`ڈbȬ�?p&�0�?6GyF�.`��?�·^B֮F�c�/�Hs8N0y��ҍ��\�I;���C�A���Ŷ�0������Y�oCհ�0� ��V�psx�"�$窚�A��.���AE������T.ْ`��"'�뤫*�=]d�l��R�U�[��WE�7����Ro��m��Y�c�rg&\����z���@Pǈjٮvt��?NM�ǜn݀�#qΖ	��ߋ[����%H]�?��M(�S('[��a��!�2�(9��ɷ|ίK�8�=�r6��J�-��z���Γ���rA(�$'�(�I�	�A�H:UK(��Evz �Is!�K��C(T+��)��C�����=�uX�
�c�b��B��g�P�
��A���>�t$�X�U2l+,�60��*|
��&�>����ð�cP֖�/��ăy�8�4�H�t#�P��1���ϵ*<<��|>O��Z���)X�40GbA, 亁���G頇�B�e��k�Q����l�e�As}7��(�MY��ʁ��ˣ�ѻ*�.��H���K��5�7�'��Z݈�A��3� \��5ĝG� |zA����C/�uҸ�����c����政}�������Li�(3�lÄ�l�Ŝj��T�����Y� �� �T��t���(�<d3L_vi��q��4����W��Ұ2]�VN}Hv��&N����s�9s�(�.L���5AF��Н1��#���%`D/���@X���L�M؎С#Q�pU9����ZIA�s-�w+�q�Yв4rHU�+��U,qg��eUaȘ�P4]��Q�u�iX��+�\�f��Q[�G$фſ����c"�R��T��\��è�����`������A0"�,-��`��C����d/l�B.��G�	�}�P�ISvŃ��/ֶ|�v�}�X̲	�o�}q�ס*Q';?N|�N�$H��g]�SϿ	�6�ZP5�L�������}����<�뮿��?����z��@�9r)�4BQ�*�`o������mGGp�I�¢�����՗_Ag������vR�#��r�(�<�EF�j����@Y�o&ׁ��*t��
*D�!�֩F�7 �nzv{���@��xf��uH��H�
���}�`��"?r�
�F��}c�-���ߗ�oB7�qH��b���J#K(W
�g��v�'���5y\u��H�~�Y�+9.tm[v�RY���"��u��!��BV��������'�����\�>'��t��畂/�49��B{��Yf��!s����r	.�gTM4�֯�$a�����#D�7s���e�!�;��5M5Q�`�E�-��Pק�(/X��*�
��Hh8�SQ$OW�,L�d;�uJI�㖥�Q�~i��@heb��;�bp�Ko�S��&)#@9���7�SmX"���5@[9o"�{�c�TD ���Q�HB���c����{�1S"��[r�`�{&=��~_��k��愾�!Ck�(jtu�ַw�'P�E֨3���<��c��@ R.�Lu��OT _,�9�&y]��|
�~G
��W��Tc�S3y`��N�������Oޙ��?x��~��s�/��ޢ��"G�	���o�|̼tЮ��E*�]FT)�:h�1R��>	A�E{[7lG�a$�����W�r�Ų"y�F8�r&�XH�A��t;�d4+%0���\���:4��^��D���Q���3�T������~\��>�x�p[%����l�hB����Q*{D؛�5d��g�1Z����U��iǱo�{n<z1yѷ����)��@$.& C�B�|���3��������� tfM!��R&�He2"_���Ơ�}������_�r"��e��5��� #����6�T�cܞ��.��d�O�0�����u��5j���?��d8�\��МzJ8���/�⊙������^%�@�#ݶ������%}�{���x乗�����H�q�bc�:L7����#�51~X_<��q������犥�#F`�q�1뮯������0H�"Ajs�^.�ݰ�x�}\����Q���R�,,N��.U<�	=s
����-�zg�-[P�DFfK���C#49��(��VV�F#ߺ
�]y"�j�p�5��։SMs�N��^&1��>	j�܌0��U8xd��z:���*��b��~���*��O�q1�!ga����#����`**ȑ"߯�>y��-�u���o��IK��r�����p�l�~����4�=Ix~""�'H���R�� �egz))nkd 0�.QՈL�(��6�l!��*�9	��(�"#�����X����;G�e�t1ޱҽ���Eĸů*�x�׃؂�PcN�g�����,v��(�Ⱥ/A�5�kA��S'Za�X�B�G�k~X$��r�get܁��(�H|ݼ�PJ�u�9�p؜i��d�u�N�F��n� &Fv !�?N��� ��<�����s��;b�}���^~�XY	�����%�7S���N�j�����%Iq뭷�.;�W�|����E	JD5B��5�* ���F_~���?�C���}��Ǒ�vۍۣ�؏/ִ��aU����6|�]��5�9&3��d��D؝]���6DMTG1�I�'���.ll�T1z�(Ç����H2&�w��"�ۅƘ�Ǎ@U�A�e��vDgG�ȡ>��K������P�}�"�0~,BQ�� �|������j}��knVxRz& R��>$ӄ~�,r�2v�F]�]-뀌��fb@M/��q~��K	�����e�ou��W#R��|=C!W�����gｍ|-)r#��
m�)Q�ؔ���X�|��ۙ���P�?� '�|2�y�]X��t<�9�֬��@(�DU=�y棧e�<y�ĭrr�j����'IA��9mܸQ~B��lhm���Jۇ��N�jX���p�Y7cu�	%�@6C��*�=�x��+0e�QȤ�"���b��~����z�I��F�6
/��.�(w[�M�T\t�d�*m�v=��B<��;�'�Q *l�ahF8����R�d�i�!O���/��/������=��2����Փ��r>#�~i�X�l�m�U��e��R"��z�̍��a�I����0�]�+�]�hD�ڥ���9�A��������'M�q�Ƣ.��0fe����T�][�3��L�D^�<8ܹ�����ß�����mq����-0= ~tG#�A���9K����	>�3+ /��H"��b�+�&�Q;+f@Y=�T�C7��B�Z8Y_�6 o����YF�*��B��p}g�Yo˲3��*+݋�_$�#iJ�!��B�?�r�Uu+�R�2sù�'�")sMA��7{2��pʜ�Y�=�6�:t-"ɏ��)r�W\-K��H,�l�<?4�    IDAT(pv<A!����9�#2�U�~��c0�r�����z:trZ��w
���XL��KNǸ�;�-D>Ӎ�N�e?��Eo �c�X���rA^;O��F,��mW�݇ _|�mZp��S�-}�es���� �Ue �B���s�r��1q@䅷����|���r=�O<��ѧ�~�q]�d��H0�)�JZ>��Y���\_��)~��-��i>�T�ʖ�a:QEŶm�㸊M�%���!����T�R��tM	����P@�nK�ʖ��5S�5�*!�dZ��(J8�`�Ϲ@um�x�!�S Q��Qv���uM��ȶf�
žN���N2F��[�5�8xqۢ�d�g��AV�t5d舤�E*C��>U!x�4�bV��6��d��#EOg��ddn#��	T� ���;������Y��KS��q��Mqܒ��Wr��0��@��V�G<�VF���V��T|�ŗ��[t�����AȔJ(��|�y������ю\.�����q�s~��'"1�J6R����_".�����~^��E��$���]*���p �P(�������E����䵟�����ڲe��@�k��@,�y�8��-��֣��p��W�K�Æ^)VI-��kf�1�
�$�m)0������G{]n����&B̷w�(%3@���C��p:+�h���-��Z�%������3�M]6K(&�QWW-��7�n��z�R�5��s�*U�\|]��7�Iv�ʄK�+���)�! ���>�J"�-&b�v�Ø�(޺�0\x���p`��UX�
mRm�4�)8b,��+��'Wc��K��k_���!<t$\�R��1s�'n¼�'X�_�vӅN�'���!����'��ۉ|�$.��}�o����"S�C	$y/�"gA��aAʙ�
).���@�^�l��4"�/'��uP�����)�y_L���φ���I,�J��v,�d�kH2�Y��Cp�"Ԓ'�rPG�*3����0�PF��|�T����\OӒ4zt�3Ba�,��═N�����l���T����*{|l~)ܮ��VbF��)f��W�2�8� "���\�3�����zћ���W���׫����C����;����N�ٮM�i46��K����Ur��^��-����;#�2o�E6�D�*���ݨ�;p�yGb���Z����w<���x�|n�d�#�����D����%L|v�I���W��-�[!��g���Uˏ���4B9,�܋9劣�,f�$DBs$s>d����ݲ+�mH�mW�2(�[����śy3��C�@臺QB�
�� �N8�^��oU�x)_���	�O�[^0E���L(�)e��މ�#�2)l���攓��ѣ`�X�|�6�AO:*��LD��A�X�L&�2��@�%��` $���IP�Y�*%!�TR�כj�
��Gf��_s>pO1����"��؁R�p�LBݔ˨p��u�d�of����}�(�{�^S�ӹ��8_O=�8�_r	L;�/ @翾�a#���F���d'��߿�Pz�O��
̛�z{�2Yse���b�RCaym�!.Sm���O�8�V,G08��9Y��;\Mu�m0���l���/��"�?����{)2|OP���X��ܭ���#L n����!L;�b{�-X� ��jdsd]�@#W"��	��%����� ��y<�x�	���G�d��c �8�q��ҒTA,D�e=��SC��^J�!հ��7���d�Xz8
G��۳	ی��O=��_��4�5Q��i<.���J$כ+�0~�'�j��EU�UB��/2���#���Ȓ∼ɯF�'�ᵿ�����^�Y\�~y3_ ��i��'�ر`d[���K�aC��>���Pf\��m��4QRV�зLͲ��Fx��Ʃ #�M���}EI�����ًˮU��r�|����&ѱ��r��q�^*t+�>�N9� 튦z͚5���/��i�C��{�C�}-�-Q��Ry̾�A�T;��Zr�����j=�6w.�o_L��-�������4�W_A�����;"��G�����_�ug��Z��0y� L;��Z׋���R0!K�����\�[�x��Ν�AA	�3i���н�;L���K=N?�6�ET�z���\%�-m<��s�~��8��q�s�t]+�_�����@u]�֌��w>�L��3�?�G����@٨E�rD;h�����R�{{0u�@�~�.x�w�ԧ?�n�8d<�\�p֦��q�ġX�� :�Au����q��? �oF��A� �Jp]P)�(Ԏ6�t��8h�-ID�~\����<��Z
�D�(:\?WAxN~��51y@�ɷO���9�������/�콉�=�����˛Ŝ��OS���#Ś>�<�%�P3��T�_ca���)�@���5~?!�-x�S�����-�y�4B!��"��(d��:���)r�vrL� $3يM�9Hi����튃C!�@ ݽI	��)�תB�ͧ��+?S�X��H�(�BX���eL�Y��ض�TO
�H�TZ�D��󨭋	�I[E��0%�L��n��Z��n2��t%μ�a�D��}ݬ�I���=�|[�w#�PC/�ɍ�g�ȭ_�7�\��$��wKPC�Bw�K�~��y�Z\t�ŒIN��-�܆��xF���*�{��iBO��b�ec�J&�u�����<��E�~��kF��aH�G�V>��x�]�י�,_�\�����=��E�;o���Gv�555����R�S���H��a?�L�p��X�VD��AȄcxh�a�I�1e���:e :��W���/����|��
���xp���
2��1����I}�eT�W!�ˠ�'���l�L2������aa$gM�5h���w$��畝0�#�4��m@�> �?��6�ۭK�$�i�_y$K���Q���_�I6���v�d�[nN�e��*z�;�~�D�ry<���@�V�O��b�"�z�"��MY'Y�)×i��8���p�3�њq�mF��_TBP,6���oi��\i��R؉��CXՄ����� �m٧sBW7�m9*�s@Xچ+�`?@�U"$�7nvc��a��Ѩ��-�b@�5�&��#��.Cѿ��s`]'���y\t�U�~�i8f߭��!=(�E���cҤ]0i�Xl��`S���'4dFkB�$������q1㎗�t�"<x�9�:�i8���3�?���������Ew����C	��)s��V�O�F���Č[?�g���&o��:��%��'l;��zz�p�Q{��_ƪ��5\t�I�nZ�M�4����Z6v��Gf"i'�7�%Dk��u!Q]%	���)�
#Ӂ;N9�n|K�E��u(��
-Ղ�N�}c*��y�E�u�Q>a��1�.�41�"�A,z�rM{7��������g�8��i��Ͼ��Χ���	GI��p�R!`�08rB��䝓'����-�[��%o��ڍk֬��U][�e�V`��Qr��(�X�J
1?o��O�K�6���ʋG�"�MNb<�Y�yxsj�ĩ`P�<���;~l���Ģ���J���P��"!lho�iuC,���d�'Pv\�Q�i0�`r������W��I�r���C��UD�u*�����^��j��ن��82٤L��]P�b�j$��JL�eC!�����ѝ�v�*,�0Bh���T�b�0����	}�l���Z��nx��!(����B�>82��hC���w*�D�<�B�b-�����_Ƃ?����D}ӳ���9�֯F��R4��r���3�k����	,�qC;�8�%�^���PB����Rl8=2��1���ZK���If����H��xjk�^ٲ���y[��]��.(�S�qO���b�۽�[��w��s&N��#X�R��D�4�z7�³��aOEצ�x�ͷp����_���Cb�h8�z�>�_�SdY�myP��l����i��IL��H����q�ᄣ��_~��o��~}ћ��BSw����ú��h��@�_���߈9o/��o8�X����}��E��-��U&���t��O�0�@-z���
�J�b�G���h����YE4��@a�QPq*��Pi��(SׄR����(��԰���JYT2x��{���7Ķ-P���6O�[��-E���������-������ר4B<|o�a��Ra��B�6ix��i��3/�G�'��<��R<1�i��U��i'a��q�rޝX[����[NB< \p�C�؝��!C������-�z�h[׋ky��� �F�gb�1�b�ɣq���auO+��1fP=���X�B5<�⧸sλ8���p�;ụ�8j��pꆠ�ҫ����u��v<9k�d z�l$bqLčW��;��>���j��Nx�����;＆���#>���:�|��n=
�v��>�Bt���2�)��#���;�){큎�6|����e�*r��ze:֮C�RO?y�{c=���6�x�(t-�B��q�����m��EuM��F�V�t�)A�\���(��5�\;��4��a4�9K^�U�Zp�	�`�c�`������+�c�Ƀ5 ?} �%L�|x���g����~��}�O?��w��dy�`�2l^�>]��	����T����|#'<��U�@Y�	��^�r�q��AG	�U����Z�����M2�?�mX��~}�����X�$��q�-�Z������֢7�����5�	S���\�(Ll������*e�\����St��X�Z�)۴���0lP?��44�Z�6��o�H<(�ش��⤖Mcۭ�F�����<�H���ۨo�Gkk7��"�jlhYU7�Ո�����}>���pߋ�c�݄��Q�G��K�w�,�d����(�nkE�]�@��7n�wͺ+W��{��C�����K�x�"�0}a.4#�>���K.�[��"�Ӆ%�/��X���U���19��MM�ش�Sr�Y|ǌ�J�8N�l��:JP�����-K��)���?/�E�O4�!���C���Y* �ʢ�:.Үpďb6�\FH㌳�����[�'�q7�N��P|.b!�����Oa�?V.[�G�} �s��}�cԍ�������0���A*r����jk<t�]_�7_t�ٱ?>��"�j����aÒo1���9\4-�5�{�D�
��^ě� ��
��gߊV�
H4I@	�O�GY��(|�*~�r�06t��>���;�
Tϔ�2|tQs�V%Q�sK¤gyWC�)Gc��#S�� �d8ܠ�<%�r�ĕJ-������|r���Y�f?�����YG�_��8��gA�����$�����	UQU��.�|�i���'AIGt�:�8�z��~p�)�b�a͘q��fH��t=�������&�uuN��69������K�:WBD+c���a��N�E�u��f�6,Ɯ+��;�a����my(��}'����특�����k;8��;���������q�5��T3���Iw:�ahA8jЋ93��'~���Y#��
f�<o�����q��~�i�w�ih[�{L�+~Y���~xr�8����XP5B�	���>5��q̾�<�n�V2l�����11\��Z���h��������E���_a�4��H:,$q��'a�1*.��3!����_��E���aT��o9�y�m~�%�g�q/�}@iI���jI��	W<��e�;6㧕JA�UΨ��l��z{�����r�ￅkA_���g_��`��V�^�ں:467c��u�%L��.�v�p�ӧ�:;d4�hnnB ��MXv�رRܸ���s��/iK�T�`�&�>C�H�c�7p ֭ۀL��ƍ��ۯA�ӔE��,)��h�9l�@z�X�r9�jkPUW���N��	�z�#���P�l�h�l;��a�=���m�}ڜ��H�n�En�+6�66����fzᆄ@B������	$�L�l��bcܛ�bɲ�h�9�̼��h��Y��Z/w-�[+�%K:s�̙�����Ƨ�.��` �&OD��	Y���pR��`{�v#�L��EP��1�|r�l`�����4T�w�����B*�b���*k
�00؊9��=?�5���l�G�������`��2���S.�^��=� (�PQU��IA�W�Ow�goÔF�o�f��6�%�<a"��nFWg+�:s���v>Y�]�O=�;�|�E|��r�ܲ��52���H+�e[�����8U����{���� �<8�}�Ĺ�4¨g E����{b��s$Pc}���hmۍ��c��߇d:���44�=H�30|�n�����Dl�X,8�<\y�f��f��*V.�3>-��MU��ܯ��9�����>��;x���P*�Ut)�H�r4aг*�l
>�E����=��&L�V��&��^x:[����Fy0���"n�_;Wl]�9����¤I&���1�ݒ�Z���hv�.�H��*�V���D�ե�6�Ld�qCa�s��.:
N6ǶX�%1P�	�h���p�ȳ�r�}0kw�s-�ͨdS`y��w���R@�p�Fd9��^�(���Ĕ���(����)�!�/7��(0:d�N�;&r�A�j
ᑻ΅�\��|�}����S��F��v;�U�q��7`Rs _��V�*q���x�����ՋS/�O���a��J���U��K�"b*X����hK�;~�nT��Ҿl/��高3�W�t�nlG��}w^9N8�k?Z�iM�r\r�]�r�A�ﶳ�z[���W(�N�R�En�gOOr��"~w�W�j����k�ak&m���\��sd*��%|��x�w�8�'�5w��b�����?��	�{:�qTCv����y�p���SŪ5kH��WO;�f�W�Y��Vn@ce�[p�Oo�G{��œ��U�)��a`�|�k8nN9��6� 1�g����1�*�.����"aP����7~G��s�7���?�M����?���-����V#P��U�\8S��Ŕ�G��(�7/���/���3�R}˺Uc~���ʦ��棛���2��s�dչ\^�ef^>����T+�Acc6n�(#�oܸQJ�MMM��3c! tuua֬Y�wn[s`�'c��;�'�����ATWע,\�l6���a����˱��_U+"Fj`XH\6#{U�Aӧa��"d ��e��8^�9M?G���PU]��hH�8}CHgr�}A��	�oチG0��@�����뙗��a���2tw�#Z"MWo�%L�y���0{�<|��_� ?���kxq�Z|��àR��}�I��qΡS��Fye��t&������w�68 ��]�)kƲ��c���tg�u>�uq�����400��G���u=���1����H&������E� ��+���-���c�b�hjlF(���.TTFD�*������Y�N��ۖ�J�X�|N=�t�رC�*�#�e�a�'�%���#�4�,:Xt�Ѩ�T����}�������'-(�mF:��?@�m���H�Dr�Vj u�>̙4�/8�	���ǿö����4h��d% �+给-���3����8i^�����~��c�k��ܶ�@zz�3�3�L�b��#e�|�^��A��SV�
��H�i��}bQ�<�G��]���t�"#��Oz}��/�(�&�����gҖL�^��y��Rc��Y����u�A�"��yc`E���=�'�TJ^l4T����ޥZP��/G�����R��7�����e�f���PuM ]daUnA��n4����A�K~��_�u�n&Y�lߺ�L�������^��D �����CM ��'�c�����q��ïa��Li���;	�i<����3%F7Q���W�c�4��;��[�1�(�/.�3    IDAT�� �`�D�4�;}�?yF�|��\�tgq�V���}��ok�b�AD�b��{��i1&���aߎ�1�8tl����+���sK��ٶ���z�h� >zw��5bl�D�r�5X��_�}��G?������/��q����^[G(V�"E�q��L`#����[	<���pϳ-x����Fj���
�D�}��8��
�񥵈VǠ�݈f_2���\�|�)F#�2�і&U����;����n�"�@���	W���d�9��Y��@.��T��N����^�lֵ�:�~�{�R}�������Owvu����%��֭;��F��~�5�K�p�����\r8�h�Lz�%�_Ϊ�*)MS<���Q8.��R�Ξ<K�4� ��ٽ�S�9O%"�5S�c`���G�y��\�S����&�x�TD)��G���iL������ 7��];����qc$�`�{衇⃕���[��
带Qx��WQYòi^J��`v⬰�CCm������84�'|�X��4�!�zڤmP�Ԍ��V��Cr��gLAE�(�v�ϠxⱿ��/��lt��	��ُl��Y�U�/Jw*���A�ð�Y��!�{��@z�l?�uw�/�@}C-�lՕ���(:�m���vt!�v�k6�8� <�q�w��M�W����� �G!�I
[����1cq����D����C8����7U9I��L�d5U5��$��Y�Ν'���W,G��.D�qDŎ����9S��	�a��Y���+1��9��?�����&䄹EU0/�w��@ȏ�� �~��{`�X�l*G��'na���T�5e֟��&�/�'��I-}+�Y�p���k�:����;���wʽB��Q��b��ٔ5�C����gc�#�������v�?�	9��܃$��Yˉ�.S"�R�@]H�R#gY�� �DI����/^�9��	k�����I"#J@�9x���B!��P�v*��M�F/�|)���y���$�q��틯Z���Nn���������/��GdeKY���@����8
TJ��2���m��p�8~u煨�5��f�o��-w�7��]���J���1�.��\~�	�b�q�1<���I�W��O:�Ϭ�}���缵���8|�<~u��8��Z|������p���ƫ�����w݉�.^���?�|�/���������룿Dn��3H"��b@'�f�g���[���~�>^ys͞��n>�^��>��h�����=��}�ƴ&��=��O9�No�W/��=y7>�
�~�}P�n��?1{�����B�����$%i��
n ��^,�����������w������Oß�Žמ����v��V����B���"ey�|�Y�AU�+:�Ӹ��EX0�&� �	�0p�C/������a{Rي_E^���Q��RXب/y����}�p�����
�>Y>㖛nZ�P[����TJ����k���/�r��[ZZP(:�}�,�DG	��3�6RjT)_�?^>�\Ĺ���m��s�ɓ'��������VV�J/?�@۞L�4�O�2~&�Ey�~�!f��jF�G X�������n������={څ���2�ಊ���\�q㥊�fv���~��HDR^u�u�1|��cLh�hyH@IԺu��d����4N�s��͘q�,%r�loÄQu���PGw2���n1uz��'��î�D��مtNG!�J��sw�2���ee�@Ѷ�IX�S��w���F�|p�I�'�Q���(B�2�Ubo��-���Gg��g�f|��������M�����ۉɓ��s~�R@����~�y�O0O�����|�QD<�Jb�{9�]��Z�,*̙3G�x˗/.E6gI�f������O��fPW�0��v=v�Z�JмY�������{�V�C��L�}eݘ�a�0��Y;7(Y@�'��Aĳ=P�>��r��<T��i'Y�!m�PE�O[�N��Ѥ�WF0��q��&1����	ç	�����C���*�}�=	hVF5N� ,X�����(�6��<�!������Ιg*�q&����+�%X������qt����d�]G���l�P&\,Fm	�ܢ3S��y��.}ˑ�L�	p3���{��{�~/�,=���h�oHq�zx	��	͌T\����}��89���*�Ġ�"�r5�c�((�q�S8r�DTEd�ò�p$�wH����at5�����p� n ���6�A�&4ajc-�4ڒ9|��s�?	��L�@��Ȍ2��Ɔ�	dRi,�ބqc�t��H璘X�Âys���]hm�Bme��9;wm���vu�A�sY�5�p;���;��k���OE�b8�[p�Egᐓ&��ݏ�S��s���{Г�<p�����b�0s�l�*Y{j�j�b�*u�ih�cgk��ƺz4�@���Jd�Q�:L�'}nմ�F�T?�^܈_,y�����p(�[P��c�SL�m
q����UpPYS�����<�_�*�$�y��4�mj6	���^���+fш`�}�X����;��"MGQ)'@����Fs�k��o@�W��,��˟��3C�l۾��2���K����Uz�t������(e�7�%)f\̲I����\N���|��$� 93;�#����
�vn���쭶CS���DyE�dT=�{d���F�	�0iB3��:::0��`�G���B&�@S�(D����r�!yQ���(�BW�|O�#���G*��^���d<��be�lk������%���X-��;0�)���Eˎ�ػ���R�`$��>�CH'���`�q��;�#_T���~��>���q��Ƣ']�e�P�~��e�s�T+*4�p��
���*?�RYY�2��#d��a�#��J�%�Ӆh�U�z���}�1�Q�s��.���$a�|�@Ww/�~g%�yCeR��lن3�>��}=�~c��q�\��	�82�&�����`�E�DJ�� 9���;�X��t�L��� �Y�-���CU�,��y�2)1�`�W�9psY(�+�0
�����q�Y�s�</��T�0PV�Ę�Q�0���ظ���(h$�80	*n����g�-�𕅑����Q}�<�:H������z~��(T�r�~�������P7�
�0�^oR� f��d�$Ar�ݡ����\)c6M�Z�}��!g��(*�Z}�F�{$9���u��'Ҭ�q8�Q�,�6�<�ʔ��Xl.��s�Ҝ�L-� <��<���/��_�r�"P�oč��9�/�2
����<3��0�tB��ie��)��NB�-M��e�d�+�Fc�r���D�eb�/�)�^ղa[i��q�EC��*,�2�E�J$d�
V�S�N�WA8\%@C�������k4�0�A���Uֈ40K�.u�Y4��hف	�f�uO'|��4I��~�(��R$�FQ��	���,��r���P�++�75��Cy����+F�����.�9D����>���ѽ����d\�A���A;�r7ŵ`SH�>�:��Ame�)�b5Gep*:tÇ����( �$�@踬��s4�jЛ�|<'����9ʨ���{t~����_s>˚Sr�6d2)EJ���&L��+WJe�@�~5��=L�P��\.+eL��+�1�\��͝;Wf�YN�"�ov�ۙ���]����=�4����̚���oBC�h����ƙb��
)�wv�!�W����4��0~,v��@2�@:����c��_^���sO�hiq�Ba]oݶY��7f��Ƈ<�]8�P8 ��r�Q���%~�d���H�^��8��:�ݹWJP�Po�.�П;���K���V����͸�nG��b#w��~dl��Ǯ��f�n ���E�)W,"G0V8����p�����P�f"�T1���r��芀���ZT����4B�	yOc �K��"@�VZn�4�����י�	�g�/"d���م�.\�K.=?�Ƀx��W�m�_�l2u8Б�L	 8{O"��h"�C�D'�F��7��*�1;�V�b:~p���>m���'���m����F�nf[vT���rN����(kc:��0P�b���$)���,8����|�v0�u[X�^D!�$�b޿t� �x|!jȄ]�y�	��LV��Y�ώ�SQ5u��%��f^paҚ�X�ҹI�n�Ɍ��v���Z�+os{f�*3���5�:��p��:Kͮ�p�X���td�[��"YC:?W`��՜Lz�Ɏ��,ɊЋw�2&7��=8����r��,>(�Tz��
_T�_QM�O�]�E��T��'p0�cfnåm�Jba��獾��}!9�T:��H�z�ur�4-'�V�s�E���ϑ>�1�� Ҷ������ݪO��O�r���_���9yj
��Jr��.R��D�f����"?	����v��C�H� N�j:'S!)&B��!w�5 �y�$m�|Nf� P�	�޽��AC�{�!?
|�mTT1��[T-���~l9������3�4X&g�Ǉ\^�pʒ����1�E���Z䔓*f,l1����@�p���
�p���W����J ��7�"ͨ��?UD�`�H�X�z���=3��-�ʘE�5��������'N{�ɧ�V][�;[l9�&YF�79��zd�sSH�p7J� O ,i�M'!�_,�2;�n7ˎ�q�mu�mg�諳d0}8蠃dޙ�[�HX �Į�-R�a�Ϊ{�mm�EG��N&=���߳���<��Jyb'�f�a�����}�8�装�չ�ӦM�̞��\��vwaT}��x�l#l۶�g̐���{�ɬ��c��e�d���������Eѓp�u�J����?G�E!P����ޡ���SU���J�V	ۦH	`s�",��{���pc���ȥ�h�Imf���:
,Yh��v؋O!Ⱥ�n#o��S�

Y� �P,����߀�D�{/.9�t\���p���ko���~��;&�9�&5�ly=z�o����@~����	'Շʲ8*���	Ȁ�~�B�abh�Ӎ����q�=⽝)��M�]���R�ᨢfG�a�,"3008�Qt���ڏ�5}8i�xl_�.V��2N9q�|8��I��d�<��Q�&��4Q`��H0�������Ü��p�M����'�P�]���"�>�{�fB$�G�s������#��g��K�s=ʜ�=���������~I��OW�e����x�{ɒܣvz�����X^'�;Wq[�*���9�·��my���k�:�#V���/σ�״�����(�\=u������3��z4@�8��*�^����K�;����x��w�zJ�/C�]sIF�t�ו�Ѳ��K�3��'��W+�^��~�'Ϸt���wܮt��=��{��)�:�^���Qz߾�����/�������K�,�{�5-�ҝ�����g�ڔ����G���~��_1��l�Q����xA���
��;C�����ߵ�<w�#��́�aT��w`oO��ј�bo��d�U�16f�Z�U	����¥>���E4���Ir7��}3` �h�Yh�z�qdY�������~(����:"3[ľ}��������~��K�!�1������P�m�/?�s� �*�R���:x]�㹔���T�f�AY�hy%�����8��tD4�ˎfLd�[8��Sq���'��w��a�������,��{џ�����k�+�g���ʲ���U���Ri8D!;�k��	hQʝ�&�i�`D�|~*�d���E�2vI�tc�jp3y)��_��)��Ԇ*<����%��7�G��Nb'N9�0��m߹eF ��|��i=��[#C:CXf_*���{?Ĥ����)R�{�0m�<��[ر7��13��ц?/�OQ���_#g��X�e^ZDw��jS��iVa"�
�����!o��!����k�?��g�G��'W��סo��\>	@�po/*�!�霋P�%�^�5�i�_9%��!R^)���SW<�A0�V�T�/(h�I�*�(Rd��"����y� �0��tOO�K��j���^�Z���B�T����\3]���'9ʁ��%�`��`��Y{���{SF�YN3o��]��Ɍv�/�O�m�2��U�jQ�A���{��!�����tI�a�S�q�^��~Ru(:�a���/��9�g��V����m=;X^��l�W}�9�X�?��L{N�R3k� @�D��$�4OMĨ�0�-T��
����dm&2.¦�b.-�^�nԎHg�V���a�EX�TD�Y��w]g�4D2��{�}/:�iEq;#7��uJ���X��4�SI�z�k��P鲽d��� 3`w��N��M"�ÈJf)R��T#���kC��( �׭�{��N
K͑�}*MjH���N`�W)��#��E����Ԣ'��a~������"BO�3�*� �K�xS0�I���W������=�{�|�%W-}�G8����!o��YZ~��	@R���#����n!���z$"�H;�s�x[N��o>�`IB�:($S�����B��f�;3ff׼y�l�Dyl��D�c@��82��Gco� �}�f����6	"�d�����s�B�l�����& �k%��ϟ��k�V�����^
J�"Q	h�NK���K��D�p8(�c��������?�K�X�ysO�`FÊ5[QD��8�4a#2N��[0:.������ؕfH�S}0T9ہ[���G�d]a���Qs��\�@E*���"��9��L�,r.�
��*�O$�+�T�W|�8\�8������Hƻ����쓏�ڏ>����(9��׍��mAo6=:{��D.�h���ߌY�
n��BL��Ǻ?�?`@A�?��!�ߖBuE&����S���;^����1�)���c��jI�,�U�����* �d.Azh7*����Sѳf-�[��N8����u���"l��G����%�$�1c�dDcuP�e~h���ݭ�Ӿձ2t��E2cH4��mO/�F��l�}�DzV<��a%������0]��N �K]w!�q������Y�y��x,6��:LW�F��Ι`�;B�nO�� ep��ٍ�J!X08�@�}V/�epį���M7Cz��lo+l�x���. /to��n���3�
R�L��f��?�`y�� a�K �t�z!��`,g���9�/ %C��f���Ixrn^`��e@ow:wi&29����2� -+
K�>*K�n^����
^�֤T����_�[p�)�"ai屝dːb���Gے@�A�<����m{�B��)����nDʂp9!�Ү�;���w(�a�����6X��c�\@�C�Ez���-C'�v4�'\hE�;Q��%z\=Mx$�����T�a�[�Ȝ:�����(A������m/������i��\�"���2�5piI�X�}�@�;P�
��v���Cc�+�^�o-������o��O��"V�Ʀ1f�dR ��^�S�h	ؾu��k�B.$_�����x�c��i�A����t'�r1 ��a�wJf��7fה%e@�&�2x`�N���b�p&L��2���y�|��5� �7!����x(�����/4�������Y��L=ϕey�<��4�5m�'S��.5���M!f�r���t�I�����!�=�^y�#�?	ˇ���҂Hm������Q ���HC�	��o��(�a  �!
�Wa���ad9�e���OQ���U�GY{������0]�tf�_z��|�4� $�9����q��)���s�4~".X|��7m[�#їD���(U���n���|�����p�`��R6��p'�m¹�B������2҃�8p�4�mB(*�������}�kb���7��{�b]g��:�2.���Ō'��H]&P(�h�b��o�#�?��Pc������	H[9���I���"�ob~�N��3���t�v������Ǎ`P$�>��-��    IDATl=�~{N8�p�߈>܀�_~�	S矆݉�X�IKȀLRP��+4̎5*���� �*�4�H��Z�)���d']�}9�>�`�D�؎`���#����r-��3+�鍲�����HF'���Hhs�mu
��{K>�ae�3�#���zcG��^ ��-p0H�df�̏�~>8l{0{'��;��϶��\뙩sM y�@f?�x=�}E!���<Pg`�G�����@�y~>裮zA�J!���Y��~X	eYh��(�h�/��-�	��� �4H��Z�q@	"iQ�,�7�{��z��|!q{�*�%�����Oא�ȣ�!c���-�A]Ȋ>�&\�^`�
��������G�-�4|�<%@	��o���*�;�OG���7�X�H�x�\�/�1PBX*(���s������
2�(�I�9zmY��sɻ��pF�U��M�)�����(�֔�V|.Ԁ.���aY�W�=����_�������ck���G7?���?f69i�զ-K2S���s�����3(	xD�!���%��Ǎ'`�7��ާ�ȢFm+V��28�%��x�q'H2K޴i��F$2���,��ez~`	�$9V��|>����a��w4x$��g4�=�%h|�Yr��:�X��ϗ,���l�F�(��VG��j��H��k����2Ҷ��O<W�Z8��{~� >ݸ��F���}	z5P�|��ZD�o¥�{*-Ҵ��/�?C:W``�i�T'���FX �ŀا��O�p�<�j�P�Dʫ>�	���Zz��2=+��L�z��߆�^y..>uN;�4�r�8��9�$;�8	T�W������p�)'`_G�|�w=�1�����Cp�8��}��cw!ѾuQ?��ɽ姉���{��w(���.n�����8<�;pҵ/�-s`��I$SD�5̂��b������߬�b����7/>�ӌ�_]�%O,CŘ�Е�E�(b��-So�b12��P�హ3�u�JXC�p����'_��'�a�$i���C.���x��gp�7oEk{/^��R~�x{� ���K�j�`�a@§ �u�)��GT0����������E��S׋h.�޼�9G"P-/�0$d��&A���F�1����L7��<M@��_��(d;��G�f-���O�8:G�R�Ն�d��B��,N�c�s]�ҷ��yd6�w�6�N��Y���+A6��b9���AЧ#O�b݄�� �yrR���X�^�T9d�O�}H�d ���qOf���(hT5saL��4�|f ��4�C�)6촗0��Ć-��e`@?l$vq:�4%�p�m�sPH�#���TC��E5��	O���6���:PX�ʧd�ֵi���l>mK;)LP�R�&\&~�U[-%i�Iw��{��)���K���S���e���d~=@�4I�X�+v�m!��H��t�$������ +]3a3peKPH�,7`P\��a<��l9�kqjnꍧ޾l��� �_=�/������ '@ؿ�[gĪk�H��j��%�M%3t�fL0+��	3�eF��m{�'��`ʿM�2E^�"3y�*K�s�r�m����p��M�}�w0s�t�!	�T+e�2+m�;��,���=��fΜ)�s�����U�;χ?���"��ϟ���H��y���c1`��d��I�J8zgP���D˱��UU5�!$��Z'�r"��{ߖ����/���qΥ�ƒG�AK�2P�++��L�� �*B�>q4֯��w����CY��wd)�0$aE ޛ�����Ӈ�B	Ԡ@�C.�V��b���e]ZP"���,BAѠ�4�f���p�����z�ɸ�;�����a䝤d"T�c�~��P6q�#��v�5Y�L�n>�q�A����ٶ��:�yV��D
'��'q�>�~��S8v�,���p�<�m	�*<#.z�gR
���K�&3�j�����(�I���.�|����9��}�[~��g!�������c7B�X����g�� R��p�u�����cO��L�¯+�ucʌ�x�ٿ����_l��\�<�:z�]��B�ͅ2��xf3�TVH���#t+YLQs#�2��H^�S2lf|�!�n+��Z���S��up�V�#�IC7hk�탽�f"[ ���3=��ܗQ7V	�?�K�*�	�X�r=h��1��d�5�G�>�J����#Q�=r����g�\,7�GJC����_��rpSC��9�8Ժ����IM�`]�m��-�ig�AEt��p���x:�qf��g��B�9^�\Z[�d��|$�2����� � �0�e@$ٺ�{O�� 1^Rm��7��Q7�D�̏�t���|z_9���� C�#��K��m��A8�����TW�3����t����z�G�)� �F���hD���)D#�f��2�@���oٚy	���L&�-���`�y��ꑔe���pI��C�"��|bd,R!����>Ӏ�#_zZ�6O�y�����`�?��_*�?�нO�z�yٜ���^y��r'�ĥ�̒1#W:�;3s�cR.��h��e,Ƕ�	�?�%�@�9o$�1�h�gƌB�#X�o,��@� �7��l]>{ڼ9y��"�	n�}�x<63t��yn|�{�e|�x#W��$)E�ܞ�ۙ����R�Յ�?�X���y,j���a��ft�z���PFf|#� �8�+�����<��1|�f3v�&P�BW\G��a�ue-јB����K�D|�fl^��X8��ne�rM�n�x�� l���Z|�y3
A�N9�݊ͭ�R�������:҉|�J��6ֵ"� ���*ʃ2c�����w/?=g{,����9}"L-���
�u��HM��+��\w��ql�c[������ Ƅ-,{�&to؎�����K/���p�'#Z���^�۔ƭw�G=���\t���xs�(�����XAt�<;�~���+}шn"�Ӌk�?	߻t4�z�c�ןWB���dڂ�Bc�Kn�'���y����p��s��soⰣNDyE�lڌX؏����6}V|�g^���jP8��������?C�a"z&
ŀ�ݲ��~��3#%����t�Y�4ݓ�Uك�9EV(<LMvM�g��;)��N>'��AuDC�Oy���ޤ�����s����TVo�� �4�Sh���F��`�������{J�u��L�;&����&aPa�� ��r�)"#��Ot��,�y��Uؾ�Ҳ��O`�
6���ɵecXسs,#�B��l \	�5O�_:�^���O�8�v��.�Tm�y(V^Z����H�c�(�ҷl�p��/`h a
_9�\������-�������2�6�>���HXyh�j	4�Lڳ���w���K���H*7$BF~��Y��H��U#���^�Sy
I�c*��"
�}���z��/D��$����t�7Jz%�����{���(�zbD�i�Ay
���]��;��a�$�R_������!7 $F���au��o]z��� �_=�/П~�7V���	ټ����9�o.�ͨ��y�n��>�R�V��k)�R7��	إ�8��	�H�"-9	���	�%�;�	�3f�O�&�s[�����f���tf�`��a �>��ҙ�˜9�ё~? ~q!�`7<(���s$�3K���$(1���L0X`�P"�3a|�����N��ރ�u´=�`��/z����G���-ht/ĐW�Q`�V�|a-�\�tnz���_y={Zp��`������I+�P��,*�Fc�죰����R,u��(��q��������8�(�w��o�G0{f�q
>�Տ��*�FE��r>��x/�L/���k�옩8��q��n�Yg-Ħ�+P]n`\�h�ϳ?�U�%�i���Il��!U,C���B�S���l/�-����3HT1n��t��v�Llڮ����Č�kp��[q�m�c���Zof;��J�j�c8�GZO��]E��l�Ef�{n��t|�&<��Wq�#/!<v6l-
#g�6Ӎ����8b^a#��^�;7���]���ZQ��f��J�al$z�x煥����/�4�]Mm�q�򛖠?X�~%[�NfGXH\�G$3Uν��56{�4��3��#Md����?��0
�"� &7���I�1�1�� j�uTG�\�O{�mt����c/�oݍ�{�`37C(TU�lLiO��JaTG8%�r��؞��6���D�DmX��	c0s|�5ԡ�"��*��Df =@w���x�;z��k����7�� �PH>n.��ǯn?G�+�ـ�qbS7��Y(��PthK+������ _1!�tl%�0�G$�(&� bҘ�"��[�p�q�Ie���`ѱGð�X��#�x�)b7JF��C�`��OQ����3���^��&��6�e�W`��sPYS�eo���O?	�6~���Nw�W�l�zQ���q�b�ko�aT��5����Ì��PS�������}�v����6���OĖݭذm�̘�m;ۤĞvt��j`���^
��>�zآ*��nN䃅�(��K�����ʉ��������$�,��?'x�2�Krb�ZC�]�� ��ymf�2q�z�,���I�R�hXDic�����-pD��Cc��^5�+��?��R����޻�rDYE%4�sȶg�Xrg6;��R�^��3ɘ{z���!PS�F4թ6�� ��̄	|�7�+y�s<3p�+��� ��N�e�� �ۋ�+��,����ϛ7O���>�L΁^f��<.���ly.*���E.'?������a�_*���<&�����vj����LN��LE�����Z��p�7��\��;o��?��n�[ր5��-�Q$�[�!vV�6�v텸������'Q�S8q�����Uؽc�+��$3��0s�L�6���;�X=�yw?��Xق`����LC�����^E�٘z��x{�.��U#�Q���F1�!7<��=��/>�<nN9�ljŷ����(X���H�K�6Z�ښ&|�~>m@դC�Ƨ��7�a��������U��5���ߊ����@o7j�����P=y2|�I���_B[{ί����&_���� f���؇XeD\���2"��r⨊���è�k�{Zp�y��Ƌfb����{�Q1�0<��hz �t���g�E��3;�Sx��?���_|1�ž�0R�>��0����H Ͽ�
N[|9��(j>d�+��p�]����@�Y��L`(�YD��Ð�ݡiErTع���=��תi�Q��GT پ�Gp�G��ڏ'�"L/�P�E4S��ee���rQ��Kkw?��?��6���A�_�6���!l�χ�Nב|>M��̮(���	��RWa�?>ه�p��c��I����3���h�3��YY�&e��νln�Z����xOt&3�o�{�8�JjFy^ݔ��w<�y�7v�K#�J�(���Ͽ�XR׽pf��0�T���+v�_x!f��~�"n������#\z�|d���x	7�p^_A�"N:v�^��`"����ڛ�O���?�¢����έ���^�wV���7���9+v|��\8=�����*q�̜�p��Xr���Қ����pɹ��x���c��#+�zS��L��;�"T�(ꏼOrVB�.��X�`WP�*L�o2*H��+(:/��|Ƞ��=��R:5?X�iQ�Z?Lҝ���p.2�l���fkh�5�3@���6Gy��&ϛrS�
���>Fؐ��M�?�����y���Ǳܫf|�����}s�;���6�`�餴iZaf���&�CJp��9fF�,�-A-���Vw���bnK��R��;��D2���P~��^�9ꨣ��M��7{�̺���zi��������&��v��iÛ�#�3�g+�T������u��qQepP�#����,��y�쩳r�,�o3V�948���Mh��B4Z	'eâ�Y��˿~9λ�����o`�'i��CX��ɂ��*(���I"ս�O_����Z,}�y����W\���_��m[�l(�@�0v<��;q+���
(�0�������]ۂ��z6֏Lg+�}�#���AS���w#��E�L =�����#��ǑS���g�?��_��5T�Eq�M����B�]pR.ƍ���-[�V|�=��.��|�d�i�$�n���G���5ԉ��N�fV�;P�?�$6l���?>v��p~���`���Q�2F���!�De+���>D#A�
A+�<���w��q�1UPs^�v���Ћo~�6�F����ל��Ok@�w�e�{��t�㊫�ƻ�~��*0e��aD}Q���L�r�����^���[Z0n�4��\~��j> �YN ��&3�*(j�|�m������t��#DiM�������C��Mh�F 9��/<_]X�1,4r�e����+>(�O�Y�J@'[9�ZTʓi��k/ ;��_<�+>���FY%�yl�1`"�OS��E�Yy��݇
��{��>��y��+��@}�[��6�4��Y�XFB]�Y\���)Zr��Y�?���I�,ۄ߿����K_q����!����~��Z<�A,V�XT���3F�ee*'m���S�\�f���M8��8��z<�����p�l�x�X�x1�4�x�=\u��X��X��c|�ګ��?�QDN�<�<<�Գ�ohġsf㏏=��O=NȄ�/}��y�(���֛���s�y���֊s/�Ͽ��L�x^��3� 4��Ǟ��9�$TĢ�����/Z�Ύv�]�g�u>X����n<�<���M��0�k�x���@(V+}rV�(O��������@$,"X2$!2�#��d�h�C�"�Hɟ�(�4�h)�K+�ە�}�	�����1��9v���>��F �%���N�w�^d�G卼1����ԝ�\��R�qv�]��7;������c�����زv��iQW� �l�hH#`M�:m�9[�� ��S�I�w�>���]�u�|�=u8��K�^E� d���=���~�i3��6*��Jnd��	�H�l��r:A��
烀L`'�����X�/��ys�� �V���|9�'	o%�Zf�����?�F�Ǆqd�t�nE��$ƌ��--�:��q�9��;�M������+� �E���a����*(E?\˅��V�d��h�o~q;>��M����Xt�\(��t;}����`_"����`��i8h�,�xW��#�+1�H����Q�1T�Ǉ0���"��������0\E��b�����E'��^�<�:~�	T����O�y������w`��!�t��J��Z���j�.BJ
��-�7s<�6����t�(l�6�M���߄��&:���g�?��x9��j�UHs�13(��e��e��H`j� ��#lcٶ.�ll�����ڇ��EB3�A�.By�#`tY��

�4�8j&��X�,����B�<vl�cqT� ��C�1Q�Mtu�`�Q�cg� Voi���>~Pua���i�(S-)g��O���
c��ɔ�`VP�&��1�I�,d��%{1�:���~>���X�+�Z32��I���-="'J#��q(�^�
5���^]ۋ{~�,:���QȪ$�)��ܰ'A����_ȤP�oł�>���1�A��*"`*�$�P�Y�*�o��{����`C��{ս�C�\s�ض�5����Q�L�!TU�l�
�A$j��.� X�e	��3���SUǳǍ°�X8e�y|E����Ig��g��&�{�bY��Y9Ɋ��S�����*%�J����B*lF�(��	v4x���<lJ?8���`�����\����?SG����$|yK���jt���(�������|2�.�s��\0�َ{o�6�x��2�E    IDAT�/�o��Wu�7�CE��L�KAҞ��^�ax�$��$ ��)0�&��g�!Y��E2�ES��:��z��k�0����#���8B2Z��H���1��Fp�Q��΀��;�w��SWF��ȵ_-f0����ݯϛ���_�~�T@��Wm���q���������/8��$uJ����k�7fl�R����/���t���f%�ff̲;3j����%v��UUٖ���dv�E���̼4VF�'��LG�f`��� �1�W9K���K�~�'�O@g �ņD;��=z�<ϑ�ű5����18`F���\Ye��px>�%�H�i�h��+;av�j��4�1�Ve����w~p���~��o���+Q3v��6Z�\��]N�و�g�(�2�	�a�}�!2�~d�Н<�|~C~���S^Q����p�,�=�V�b�pzY5������M�6����y.�!��Y6T3�XU�T�L_~Xp�6��s��Kǯ}K�}��F�P��>SE8����WTX���g����N:���r��A)Z�E�Vc��Q������=���G߀�tءf��y���E�h!-�������Hy�q;L�s�� �P�����]G�B��!����M�O�-+��O�P�K �d%ӫ��E��]�zU��"W����eHZ�*ꑰ\��i�?�kG�_��<�DN=d,&k���p���8v�xiS/6쳡���k�QT���g�=n ���]8m��t�"L�� �_b0�Y��"�!�I�,���&M{�>p4�jm"�xcE��g�?G��
�_��,p�O���-=�Mrb2��:o��o�/��;J��Z��uwuN�G9KI ��9�1��d��s4L6��$�Adl�19BB9�4y�s��~ޞ���{�պk}��֌�����k�y��O����e�2y07��ue�9J�|�o�XN�Vl�(�-��S)�����/C-�D2eX���H~)2���
���+��R�䊸CQ���i��]�
�[׾�rH�Nd>æÚ�}�q�]�[�����z�Dō+,��(�;@��%UrP(p��f*w��%g�3���>�p�sӛ�b$�qS*f)�&\(&�|]#i�f�	)e����k����#h�z�ZT�>�
���_-tI��)�r���O"'h9�b���z�m8o֮�}m%/��!��W��x"K��ل��o�*z�|�eP%�V�b�F�
ͫ�����3��d�y���#��Շ��Gۙ"j`����g�L$Кl�꘧���|N3�Aio�*Y��\����Nܘ@������x��_~�p�(�D�*U���V���y�G�n\�B~#?K�����6p��FrS;E Y�C�5�����9�N��V��uvt��I�jZȞ�>��M6'Ҟ���{׈wZ���V�\��TMk��y�*u�7������n@���`���fQ�����2���B�|u.t,u)|n�	�hlj�����[na~�F����X��L2ŉ�Ƕ;����}E���7>�
!㌰�;O���u�rxȧs��Eʒ�`L]}�X�&b��L�E���=cC)�x��#��7�%_RNw�HE��,���q-˸d�55粘	�͈QCi�褐*�5��J�u���k�ܟ�g��j_N �?F������3*Dl+_C�W���g��l�JJ�"44�.r��Ǡq����o�s����	�ɒդ�0TQ��}�I
��\�LCc�v��9,Gg��&����ł�$%�*��ԓ��3���WJN�M�2��5x��T��i|�U��RN��!�Y�:��#g��&,%W��获C��g��ڕ����fШ1t�Y�me_�%ɺ����31���OD3��l?��;/ڏAnp�Sd�}�VVF-
O��(+\9��=.�OW�']H�>��9J���Ɔ������i����ҙ�+o{��Vv���Y�@��H4�O������q��=i�@.Ս��"��Q�;���]ɘ8M�W������^������s
�Q__P�i�q��Xu���.��c,�+SiM_�B�X&�qPH'�,4�(y�U�J��9���g���t������}���M���ƴ�㔼/O!�a��q,o��K%\Zp�l^�\�K�P"�+�2@-�\�,��������$#�W/���.a�Q2�rѦ�Q�d���y�F�>��Uu�Q�F�-@WZ��N�!b�^�.���@�3�ӧ���:}k�%���3�ZGЗ-`�T �c㯂��u@�^�����Hbto�=	���w@�׽��*Q����L�d�K��W��Xs-2UM��?06�q|�1D2��y�yT��r��[��?�����S��1��Q��?^��{��tʘq��n}�n���5ٖ�KuC�t���[���	�Wg��tvv��AtU���n>2wp֜�T��C���:^gO��|k�/Y��U���J{ٲe�k5��YU���U ���zм��8��Qh�]�u�ϴ0���uZl�� Y���s�O����hѡ6�f�Z8D�Z���O�|�J�Z������U�>��+3gΤ;W`��Oe��O2l�4|�����%X�F\?e��!+�+�*{L`H.���2���^�����#˘�[���(���a!�ט�x"���'pHW*弢a}fv��x�~��Л��͐�������]�	2��vFו�}�"A�{}�8��i����_�,=i��]�����H۶Ɍ������)�RDBj���G��\�����I��ͻ��b ������S`��N�2t.^M[w�h�ab�4�9��k��J��|_)�֣��lx3�ͪ�[�KΊ���ts��yoo��3�������g��ʃ��M_������p�����ky��ad*6����>S5�������q�ө�Ză����ɛs�Ig�EW��WuS,��aJ�+�<�;ױ�fn<�WlGJ��4�h�ެdQ��x�w�~�J�\���T��4�[o��8��ݦOf��z�%5��R�z�wVp{�$sN*���w�v�=o���n�HE�M��Aq�r��uK.>~��e�	=��A�rۢ,U�g�6���W�c}{����(������C�a���� ���i�Q)U�N/�`�.���s�`y�K>�d��l�,39�H�`�E����`���s�o��c��h[Iw:���,YW��R����3x��
J�����ߑ4��A�
8����=�@���VW@��5�7u��M��.��4�Y[%��X�ׅ�Ib�)�����J�/�{�r*�? �"�pfӔ;;	�=8�n��:��sX�(��F2J�+f	�)J��8t�m��]�|	̸�|#7�i$%�w��bՒU��]~�*\j��@�/�>�R�N�b��Qo��Zs�֪n�f0��8���`������(r�$~���J2�>��J�{g�P$�ЛW�b�H�ir��>x�aS9�!�?�ب��ǳO�X���Z��l2���RUgPTK{՚����um�Ñ��ES��}Ӣև��B��4�-2@���"�6j�k;�N-m���Q#�<J��/@��]N ��x��Ș*Cձ����ݝ��׌[�m�oU�:��7A��i��Xj�릒H'�yj_j��{c�1 w�6"�i����J׹�=�]���`�Y���b���yUsc3	Y̺<���[9���9�S��n�t�#?�ou`�������RDf����|�u�P�by�rJs�'m��kFv:M 5v�N�6��x�+;]�����g�d����r�����A)� ���L�c��Ǚ�eb �]7�'kv���e�u�q9�7F�q2Ke4�k�T��p�t%C������u�-��h�8�+	�+U�g g���5k9��_s�E���?r��ғ)p�)�Ү�%�L�d���h�]���$�QN���i�3�l~3��7�z�%��p�����n��oVb�Z(���N��$�:�t���n����
��a>��k��yЌy��;	�ܜv���l�<��g�u��4�| �@݀�[��E.��l��&��Ã��V��i�n���]+��՝e��jQ�!�d���53�`��!�v;�e��
Xd]A��0myx���x�O���$�m��`��]�hT��s����n
��u<�\����*��"RŁ��fCf\�
?v�B!�+������-	�7&��	P��z=�I��t`�����7l��IW��▶�� �JY���^�v�ʩ��H�c�����N��RF��d��]��ث�<��!�W�I'	H.wW٦Ի�Y���Y���e�p6u�&Q.�p�YF772sƯx��U���W�a#�Rt��%�*�ԇ�x�̞�{p�3�A�pR��B��-NΟu$���p냏S4���ZS!��W��pW�,����Nf���=�$��dKQ��0�L�`%�_��3~��n3�L|3硯 O��Ͻ���ꆌ �H��Z6�T7SF�c���g�1�����M�B�����?�}�U�f{��H�~i8Sա�b��f � }�j���H�_6i��"V���֯@Y�G�����p��!7��.�?i��~+Ȫ��r b:�[ԕ�w9}�V������|c��/�ydw{g_�?1���ڶ?U�ĵm�L����)�X��O�l&O�T6� K&����e�@]_�c}��k���l��ـ� _��:Ĵ��o������~�Z����
]+=�I����Y����k�6�H�ڗ^��ՂW�r�ut^p�V݈���%�ԶڢE�~8&��z�������ͭid�����E?�����﾿��SOc�cO��3.$�<���C���ˁ�M�YAa9�B�b����..,g����YH�1sՒ�bQ��Ր��ɬD�Z(�Ep�tJ�^S*�}�𺌯u�������=��>|�鄘�����<q�LFr��Q��O4�0֕!�]����pz�eH}d���HZ	�G7�*=��Ic��?���a^���!���}E�[��f�JN>l?n<w^~�^��K*M����ڴM����&��=޺j���@���L��v���`�{���p�=�X6��h��p!��~��*���1�)H�g��8�����C��%Za���y�a�AB>�	ڙ��#�	�� /��?=�*vx�&�.9�AS���4�U �-�(���%]�x�MO���-��; ���L7����-�X��;��:E%[���>^���;�|�u)�p#��F4eR"_��ƪT2:%�y�׿��l9����?�&��"�Lֻ�*�\��E�z\z�ct'3l��xn�ho|��{IR�ɜ�~�Y�:�m����֥(D�FHW��6���}���)�Ur�M�og|���W�ʨ(829�~'�d�0�mw����.��m^��g��bI���U����e�P9Oc��A�,�1��~\���r؁f�<�R���n��0�x?��<C!:�/d�ĭ˧
����M��S�D,�^�0��PB����9k�I\p�&������Wc�@L�|~��X.
�uv����-+W�iw�������X�S[�Q�lé�M��꫐�k��47v��l����gQG
�C�B��*R�_�ug���a޻k����p��NL�ƿ��3���6np��ٟ���
�]F4R
h�o��N�0�x��&`��������H��.좉�1��Q2�b��9s�j�X$=+W W�`��\,�yI��G�����ö���`����7~w^}������T�`�P@'	��T�2�j�x�n�X�vTmTM��T����H�sjwE,���f>��������-@V%,P����Z�[��kj>�z^t��/@����"A-|������f PV{^��Y�M�S���̓���9�0����[�4F��E�T'A���gٌBf���D>C{�zZ����r�c�}��4p�����ߝ�f�����܊+:�����]er7nw	��LY9�J�*�s:h�rI���-�D�f
y�0�Bգ�RH	)杔<nҥ�i5�X�HL+�d����e�h�����ؖ���Ȓ~dي%�|�y\��9�:��8|$�uqG�q
;h��z�A������O�(:��/Г��_ibC��B0�բc�Hu�L�68��sߓ�7���kI�&N��o�œ/��;�%�mk��w���NӸ���X�ә	�U����^6v&?��"�>�"�Ʒ�Ϙ ��yk~�Q���҈-y{AIW3N��s�Cn-)����O��d�;��э|��?���K��6����g��?�ɴ��g}%�\q�_H�((I- ���!\%7e��ic�$c��YIkNS'�m���(���_L0ڝ��Kf�U�W��Y0��y�(�����"n�ҡa�Eȓq��k-�Pr�z�J�Q�������]��I������,��+�.�x� Zr�����2���檋�b���I����[5�	E�����������=h$I�t�"+"��p��e��/�u9�d#6��P�_�P_���KOb�QJL����R�P&�M[����01o3�;DږәIʸ�yf� [���/|��<�����Y*�t������}s5��6����JU���e���)�~)�&u%���6��8���IG�#gl�m7�KO�G�G,m��o~�UY7�z?9GA�������X�����Uy��k}�&��	
]��t�<i2����_��%�H�-�%y���j�(f�?{n�gY'��ǻ���'�T�aQJt3*����w��/����ˊM��s-�)�93��	�NP3@�%����s��7�Oa�F��p�*��4���ʦ������%|�o�d���Ē���)Ű������ݷ��}mki���;x,?����+G����υ/�����t�^��ۿnԖ��>�k��ͅbـ��S�4U�����K5��[`�r����ل��՛6x��U`(�P����4�L.pj���/`�&]�_����о�g�C`�}�Z����`����G��<5��6b��u�jA�����E�ޟi��	t�W3�k�8:�*~m#��S+^mz�V�W�In��=1���N���A�})��UY��;��;����GFLږs3�c�ґ�xC�?B8h�ϦL���_�$3|���2��X�r�HأA�ɸ1q�ݔr1�:屢f�_	�.D������I��R��f�&W?�z	K>����f��^��Og����_�.S[8���4a�i���C��������I6t������,���X���	t�t�JC(��nƯ�K�k-C��?]!���g�ϙ�����ư�&nn��l��|�.��D��s���}T�%*�fyr��JmA���D�yv[O�})�d��Mdq�bY��K�!��c�2I�p8
x��4����/?8Ȑ�QƍŤ��ȣD��6���ZH�0��;߯��&�dن�FI!)��-�2����T;�h�m����D��Ǘ�d�ޛp�ө������*��ॏVp�ܗ���nCR��J�Rt�n�5����,��]�3%ӱ���QH)d�����N`�ibg	Z6���5�_���u3bx����%����ʞӶ,�z�s��v�D
�(y
��$�����-a��1�_�������CHNub����� ם{�9(�c��x%������{��ӵI��:2%���l��8~��L�zKn�V&����D�r� �n�<��yks^~��ɕy��ͣ$C� =R�����#�I��'a���k��]+��v?V���ISG����~�5��M$UV{e�!`E��,绹3Y�,�q��I��J=L�2���0>ZT����3��Y?�!#�;����1���ۻ��������9t�l?��Mn�d��(�_��W�w�Jª�vɫ��]0-v��lYksoS�x�W�w~�ڵ`���Y��,���s��H�؃�U��,��E�@BF�?��\�y�i������;<����qg��#h�Bw9@��w�>��<��n��?칙{���Q�n��nT@�OW,���E�S��8f�]����DSy�}A|U��M���x��L)l5��/[:zM͂UI��E.n�G��.Pl`�    IDAT���C���"�i�W����\_ں����j�Z\�t�:ǚ4��׹Ԍhj5��M��5�^�qt��]衅��ׂF��r�-��N�}�s,EKKcF�fC�Z֭o���54ұa=�`���#{�W\{#&o͙W�` �=eёT���b� �Gp������8�������P��&����}^\jq'zF�f�n9B8-�b/��0�TG%˨	����#�/}�ϸ���6SFF��OG1��9�e�<4��m6��s*7]w+SF5r�9�p�!�2q���n`䨡�:b��\�����,��W��r�%�2���ߵ��b��Λ��J��EI�8E��G���7���d�9/���?�f�铸��x�{|���tǮ���$�:��Z�^7�����ܞ �|�ր��zA����8�9%}�\.b�3F����U�H*�+��}!��e\��s8��C��O�y�]Y��B���S�u����BC�ބ�UO������/l1�e�&I��>�G�%W��%�pQ��v8	�W��UG��h�TGQ֨��F�n=\|ۣ��s�hA�X!��"�n����j"O�EJ�@���~�u���b=.$����k�����4L�[	b~REyo�ˤ�UHJ��s�q��/ɝ/~N62W�`z�y�dL�}%c��0�ؑziԋ%�����~=o=�`5��Ӥ�-��ݧr�ow��]2A@�M6c�2�����f����Y1�s�|��&�`�)�x���]����MI�?�*{�=�8��
��6y�oƎ8��n���X���I1���2]q0mIN�����d��5���`.>qO�z�M����{�������冡��t� �������X�4�Iw�N�7����k8��m9d�M�y�[|�`��Q�{^��2,Ye���^�`R��]8M�~}�����	�'OP�/�٠w_�#����/Ip�f��Q[T��2����^�j5^��8��j3W7z�����l-�E?7���/f-�9��~%�Ȕm<��r��bꦣM�1_*����J����9��(�/hHt.W+��1[����#���ё��y�_�s�G�xn3 l*O=D�L�aj�K��JT���W}��l:��WOgP���MW�. U��^����yN�
�T���o�����~��hj�J[�i�.��@Z`�s���q�f���Z|h;_ �sS�]���?��c���O���i��t:��W�'p8�����nZ�h�*ܜߪuL�0�AM�tv�ٟ
�X�r;l����J��sO���Fm�-�_r-�����!V��آ-@��E*K�b�)c	�}��QB�:����T܍-?C�q�*9�x-���5C/��g���q��D��&�i�I�J�;H'J8�"~�rC�ClX��R!͎�Lf�}��n�s.a���p��N�ⳏeʤa4m4�A�$�ߋ]�3n���(���i��&M*2oC����+'yv��TVϦ��I���$b��!ss�\x����'��ŗ�e�q�a�L�;�5�%l�m�ӘX��p g1�]�P(�qjn�c:�]�yE�� +@Կ�:���t���d{�4ZX��ݖM��!ӟ�t_�G�j�~�~_~��.�D�C=���=�A��&�l�ӯ��o}Bd�4�rn<������ P��L�D�u%���F[&��|�s""Y.\�$�5Ux��C�S��.��w���{^� ��M��������5]�������T���%2�N�G��Ma�
U�y���'�{��Gm{w��f�q��fU�rE�Z~o��~�e*)��l�j�Z�'LR�7c�Q<r��z��4����s��Q��̕�eI0s��^#�r����sa�͆�P@������ba�<�ʍH�ȧT �d�<x���o}�O۲�%-�|E �p��v�ǐ
�_y(����G^~�Rx�t��$�t:|FB̧٤���+��#��[^&er֝����a��+y�3>��3��<n�Ӯ����$�+~:M(������UN��k$�-Ƈ����ͻ�f�^N��Y��������RᩐVN�â� �z]~$;L����>���WS���̖h��Թ�M�k��=x���M����D���/��[���S�>P�ט���/dm�u=��2��͒�C�K��LN}�`�j9V��@$nŉCr_1�+E�Lr\cc=ݱ>*/�h����^e%yݸ
q��5}�>w<���MLݨ/ۨ�~륧喬l�*���Y\�!wtwU=͛����5�V���X�����W���^�vU�eU�f�L�j\��^�B��(�8�u��tk-�tL�p�\�K�c	�����?�xs<Y����F�Y,�j^�v-�M@,��kE���d3[�7���fs��XI���_S��h]�P�m�oe� �
uL�^>����W���>��������ӹ�{�5�Rd�~��A�
/$J��>Êٜ��O"ٹ�w�|�d*���H�4 hE�dd����߁�ncê����4�lYvʭ�[#Ih�I�
zh�4�ɸ��Ļ��v��Y�����r�s��G���9�����q���p�'s��;b�9:֭1���%/4�4��o|�O{ZX��o�����q�ŧ2�g�z��z���r�a�:{��cާ̛�6{O��ͷ��qW�����nR-e!\�>r	�e�Op�I$�ZAS�(��,�o���PV	!������!Z���4�ymΕ�R`p�ŷ�}���ʘ�cM4p}}#��+ӧM'S�w����;�{[p�[��=�4�K�\�I��E�ԥ�V�T�lE�o�8=�9vvs�>�p��� �ƫ����Y�tp��X�����E��(�K�Mƶ��ɭw�rF����ɛ���S��H���
u>���~���8�����<�%�6��&
U�e ��<�]�0��0�2>rY�|��Qw�c=8r�l?*ċW�+]��wq�3���W@�x2���:�2`q:	T�Xݫ8c�	\pԎX�B�rV�� ��\� �*-�}�$�9�ŵ��u�M�2ao��#V��-�y(B��"�mg�!En��8�{���/�O)�B��2�t�e�e�B(�K1)j3��_��3�I7�J:8
ٗ�k���HΝ�3���������Nb�]'����y�}C'�F���_����Ek�t�k�9��.�hr1��y��/�|���c�iS0�R��e�$�:}�>ܽk��W�s��S��I/7�}װItg���7��%�ٞC������T��1���@ؾs}%�UcS.�*� �	�����/5�o��I5y���%9��Tؗ�8JJ�s�kT�EO&�2]4D��3��Ƅ�,� ��^��E�3Ge�����C�|Ė�7*:�7�Q����wŬ�A�T1ͳU�
����Fţ�E��� W�W�@���V��UI����}���6�lcZ��jU��l&`(��&��U�$+��Z�[�s��kd7-2�?}U���O>�)�U�Xk��c��Z=jUx-�M����X���uz���N�ln%��{�viu���EU��p����9ʴ���������.��j������r�1�pɕ�0y۽����W��]vӖ-џuR�sPW?�Bw�|�2�z��E#v�z.��F�ǩg^�W�ʃ�=��!B(�@�;��;Lg�K���[/�t��8�X����z8�k�W��۝rmD:���J׸�p��o���~�C>�C~wk�K�hs�q����=�/<�df��M�H�ۦ9�&��S,籂~�u���O���
���Gg���ѭ�_����2�hChgd�O]��d?�t?M� �"<������O�a�1��2�Lf^�_���{�Q���0�d��閝>���"��p��N,ځ\qY|�=�*��X�.��R&���������T��c�����M�ճb�b~�a�8.�C뭷�W|,�wq��Hz%��h\L]�̕�-����j��	)H5�1�fuT����.��,������U� ��{8��yZ�S��!�,^;æ#�;ʔ26n�>.`S�"U�Á������t�Jd�a�b<;K4yˤ�}����GoG)�ëy7%�����O~��ۼ���(C�i�|�ڱK��J�o�cTS�\��Ƀ��4cw*"'z�<���<��2�#I�J,X�fP��ҹ�4�l���+O�Փ7r��#h��Y/\0����4M�~$�J�@��xo�3�ߟ�?��7?��xh8Ew�d�y��I(���
�~������
Q��9�M^h�h�����j�:Ҝp˫���);m��*fm?�sf��#o���g�I#9k�Il6f\�4���b5��Y(��[�g�ǂ�=�t��Ĭf��
o9��N�ȓ/}�U��4�, ���U�:��9-B�kG��㺳wgq�|�m؃&�1�����`�C�ۛg��1K��ĽaCH����U�	����G@�_�j ��W�U�:ϚaX̀F�n"�M�����s2��?����>����ͧ Ĳ�/\^b���PH��)��X��;N=궃&?���Ս���
�ן��p�
W�a,[V�v��V�%?�Lj?L�ZūZ|�W�~��k�_V�Ud-,E`(���\!oZ�I�[��U���$�U�,��q򺰴���6����-��ѫ�V���77�|� ��]��Uk�����ր_�[s��y�up�:�v����U]6-�ѣG������z{?z�_v	Guǝ<���7��+��Kڴ�
�!�B�\,Kk]�E̹y&��}�l?�����2un����񏄢�����s�!��_�h��i+��źn8��g��3I)R4���@�L
e|��[��.���9g��?�\�7K�x������+�:4�9g��n��M�w_��hmm��IIhn>��[�z��÷��%�y7����=��8���{R�8�;�l!EG�:�w����ӟ������e+7]43.z�����-�L�3�뎌M*���ظ�A|���>p�������%�%D�Ҍۘ�T��3X�<�:��wcw�0�!Lp�9��{�X��"C�\��Ƣ%�yi�'x['��'�k�LA��~�z�ϕa���bU墊[��Ί���ᢥ�E��[�;�ٲ�p�H��'_�ә���Ƭ;^�5x�rW�&R���s�	�S7�7��a�U�����������׾^BZQ���L��	
4:�����al�l*���1ݖ|!O:��W��[�tq�ms)�؊vi�Cn�b7N�w��p�	!e�D��d:%�P�1����KSp��O���L� �������-g1�A�D�B�kBldu?��y轕��G����R`���p�N|����)��fr���PT�]��kD��.9�{_k㡗?��oAx�qUסbil�l�I��\�k�6�9�V�PlWw�jfm?�sf��#o����o�<x����)|�m����0�N��*�y�$�\���s�"�k��3c����<��r�ۋ)�L W�f�;�!*��@�I��v]�տۏ���)ݔ�L�8H6X%Z����ִŋ���BӁ0�/��U����5��gNq�����/+�Z�n4�U���|_Ӹ�����S�@'���X�ހ�����
w�J�gD.�RD��ٕ̪
2�)U�2�>�5K9x��39j����ި�~��g��Y�V{���p���� Pms��m���P���
�
��ꪬ�!M3nm�9�>���[`. 5G��V�Wk�����u1iq�U��#V�-�7پ�V��,l��Vf?��	|uN�M���_�ՂA� ]���H@������Ӡ���\�U�v��a��4 )�˜�T���+��gOf�v*�{,��~6�v������E�_�A��H"��S��Oź�x��k�y����~��!<M��W��O�s�=5�l��Y~}��噇�+^<r�6���kK�v��|��w��T1C]�Pb�4�lC.Z]1���1��X�w��ɤ�|����ϻ�K.����ʯ�;o�v�m'�>f?�-��O?y����`	��a�C��N�X��!�m���w*�9��۰���,��#::V3t���
���a��,�����T��Oۏ�wیs��c�pEw�K�j"�2�p��f��Y>�H):)�Pp�&*[�C�7DQ�)uJuSq����\&�-��+��W�lL���ؒ�����.�m�-�6�᭿Ȃ��|�&F7Q���� R'��[�"Ѥ1ϛ�-��RW)N�Q�N:����u'Q��[.9�=�z�㽄�^z�I��<��
�{��x�M��(QN��'��d���4�>���\NTu��"5�+b�Ժtq��/���B
�-��1�}X���*���g�S�Ү��|~�7i�š���z���`��_��X���H|w��+��z�L�@@��~��(,i@��"�p��sn|����"#H��9���3o�yLo�R:nx$Ҳ[�&5���������t+�%��i�G�d�::rrM�ɕ��.�]UG�u����]v����^|�BCvŉ�YF�i�ߘ�r&G���ʃX�!͉��'J�*b��r�y����ז��oA�H�ky��Yl3��G���~C%:w��o:�/�d�##D�s�;d/.�o(s�����.��4��	O�?�1��ة\�S;����W��ߟ@{
�=�n���ɸC��^J�v�ĵgmϚ2�u��J\���k�\t�M��/��"�'����	�l��*u3����"e�c��^�|V�ǌ����(ꊮMc�k�`��TLW�'�@��`n��P&�7RG�R�����[��l�Sn�/b�F�|����X��KZ%I��K�� ���w�S��D��}���Y�����\ZD͒p]�e�!�\���@Q��j��t�ڮ��� ��e���N�����BVT�k_:��:�^��U��9U뵙�&���oU��uA�Hv&���1��{�@�����^�/@Ǯ��ҹ,S7�nX�}==|^��9g=¡ {�3{�i�����d�.\w�C����wEY���"�r㩸it{ذ�|���L��[���}�0|��?�(.��&n�}�-uF��+9�x`Ν�:���P�,Y���Kb}1DV.�2�$�d�������U`tȉe۬i�%���>`������sn��"}�^�t�vX��l�ϿYNG�^���k��C�{��s���H.M�k=#�eN9dv�z4;i�d�uM��ꇼ��t��9�Ys���7^�|)����7��.P��@>W2���m
�^*���u�w��*&���-�XM����+�*J�#�P"�\�'�����7;N`�m&�����c�1m��H%3��pݵײ�S����y�K�[�E�q4iU�~i�-JꙖ-�~?�l�d������6n0�Zq8,��a-�V��]�q�%�c�)Q��~�>)�X�f��h1=�!�L�T���xq��i28q:>�����o���6p7���Տ�3���|���Ksu����˃�c1W>�S����$�]sRG�"�\=���h�����]�J&t`g�)Ǹ����or���JS���6NWؼ��l��%	�x��,�7����.B�P���>�M���')V|�5�uß�}ğ^]�s�d2�2�L�m�\0s�Z��3o~��b��K��j��<X}�9@�ǋ��W���+�Y����BQ�LJZ���C|̽�@ֵ�9��y�����'����Y�݉G_\�}��Fi�8R�8�%��}=]"�=Ȣb��0,x�d,IpΣ��^�RN�3�ݸ��a<������R���	�(qVv�ҵ遂;A(��Cy����Y��#λψ	���Q��$ᾕ��4֤
|�j=y���̤ͫ�^�On����Z�5{X37�(?�$�����{��}����5�2���]RV����s�('9�"���z�U�w|Ug�\!t8�s��%*���`����Y|�k9|�a��9|��6
J��Q��ߟ��f�"�V��l� ��M��e���t��T5ZT`%@2x��p-�q�!�	Xk@(�W��J\ճ>p��kmq��_�5��ɮU�o0������$    IDAT��Y��:��<k.��db#ֺ�hU�5C��]�c��hq���~j6�5ɚo��}��P�BD;�U��w�ר�����K�Lu��~Jt�������8��8��c�u�����+�=u\3���AFG�������ę)�-����2v�����yϱ�^�p�A�qѹ����P����qcy���X��G�~�mƍ�&�ǚ
�ڇޢ���������T"A!�1�cXK��8�+������]wۻ<���8\6R���a\t����ɛ��KiNgJ.wu&6]t�-ʣ�B�T$2|�	�(���%}j7eEu��xMJ[���$��w�:�g^��{�x��-Y�S0�z�1wd��ԑ��#�fNm��p�c�O��e\ьV[1��wŁL�*��
�l��y�s	g�k	��+/1c�"�zcb	�1硇�y�i������w��.gV]E͖�D��ˀ�©�h!�к�[3Lh	��cO�kd��������E���K9v�f����sƎ��7���+���HGG�EX)�!�/�����o3����t���b��I�<�^��<��|�|=I�G����-L���`�\u�1{Q���{.[5��=�����s�y��&���Z���k(�9s�-�|pЌU��㖛�jS�х+:X�b�c6���.�����iGȘ���=l�r�E�3�oS�|٢7m�[���W�� N�a��M��c�Aa�8s'��g'�{�XpEo�YȨHw����6�ŭW�_����/�A�aٜM�m�,�lفG�(v���^{4֧9������$�(t,��&p��;�������dF�0��hO���ܑ���so��_�� �7��wKb�q߫���8s9��b7�:�'_��?��/
�#�dm\�x�.Y�0�T����r���\:�@^^W����`�ʺ��:�c���ޏ�~�����;bBw����\,�R`� Hk�m�楪�O�s�i�����m�IWU���O�kmu=_qa�]�u�v�T�x6!?��\r��A���M�osծ���Q��+k�b�INQ�n�	�p�*�+)±��8<���'�y�_��o�Q��Kf�-Y�)�ͪ\6s�iӦ�r���0�{�	UŪ���NU�in��e�VU��%@U����?՜^�iV/p־�@m��_��s�9iQ ��"A7/�k�P����1��n�9o}գ�8���M���@VE��[-ze��ZI�FswK��9��_ӵ�j�U���}g�S1<�J����ж�}�ڝ]vޑ}�ُ'�{gd0��a��#i�8��*��M��4��n���jt��w[Kc�L�R>��� �s2zp�tr�:��%l��%_(j<���~r%yw3�R��젮��d*N&�0�<����=�L�65눣8���㸹d�.��~F��s��φ��<����$?�ɻJ��6˃' �?�X�u��+���/a勔����oV���B_>���v�}'q�c����4��B��K<W�YԍX�<��0�r�R6e4�ᠤoN��Q��ƕ� ]�a��@�p>��U%��h�����PN�QW���w�c ��5�2r�(3�^�a'�2��kS�O[$��y��mE���t�VЈ��S���)���)�cց#p�:��s;q
��;�:�����s$��3��#an�2��xC|�:�)��L�>;�mN�2xI��(�SH�q[aӪ�$��?���!�Q��~T2�,A���3U�c7��� D�9���T��,�d�Yr����7�u�k�7�sN�<Ow����MX^��Nv�2�'�:���z�������g�h�2t	�H;�)���i#ן�;��때��w�[�.{���&���R���a�X,W�E�:hw5�R0��o���b�����}yh�j��u��#M�A5!t )Ͷ�V2l�O\�+�-�cƟ擊�1��l�B.�ug��=�����|�t� #9��ǻx��7ν�]>��S�x�*��q��/���m{�u��5;���k�����6W ��#�D���N�A�?��c!��=G�?���X��ޡn�TEe�g�9c�����-x�2�?���`l�:�4`)})5�V"����V>�

U�YG�4�Zm�WcW��%1Τ��Q�^�nP�0�K�Q���>Mӽ�ʪ��W9N'��m�1z�\,S����XLjE�/�y��]�4DYְ�Y�:q�����sl�/���)�ב���7�W6|������]}N�/d�TհLU���M�U���@~��P���,_��0�Pn����G��}4��=�cc�i�Lo��BH(�@HN='@B�@5B
��z���n3OW/{o�����;�u�=��wÝ���cI{Kci�[,����!j��u��Zߵcof���7#T��7ݯI$�﬩WW��7b��o>N#�f�
�l>g@�)�S���/P`k����թ�vSoZ=� ����)�p��y<n�Q*F$k�.^���z\*�f���[�ڼ�l�`�?�sK�,��9��w[�����o�?�`���}�axH��?�IQ*��u�V�聋�!"���	Z!?��hС<�K:�����Ƨ�}�9?���Q�2��ok��G�[~\_���\eu{�ڕ2�S�\$���q���r�=�G��p����]O�I��PX��g�vsv�&:�Aj�M|g�4z���}P�*R�(�cs���QMō��*{qo6�}���s�-&/�N��z8FvD����`�D{��S0{[\/�H�@����0�j�G\�0�I4�Ic?j�uGLnu`e��5�����_���դ�Y���C9�{'zw�F�����q����IM�2j�1���G�P�@؃����E��l�Z�g��9�V�巗����S8��E|�j-o�5�����m��D��ٚ&*bs�$���:O~�C�},#f1h��7��U<Xn�m��Yuc��7�jn#�H#�X$@�Z�;���NܗcL"�F�\2��`$D��3�Pc��Ql�K����s���5�z f�S�l�x��j�@�
�$������Bo}b�<�	n�d2�,�T��.��H"x6,�7�هcL�kW��%�'d}�?�7أf3H�x�[����v;̀�_����n5�*2�IX^�ý��q㥇p��k��?�c0:�J �#"�@-#`�pGz�uj��۞<��j�����c㍌�ۻ�s���I��禧�qݣ���0�\�!�S۰��'��������ҟ��_~���C|�ڇ��Aț�����kd��*?��A�H�z"�\�h�R��O��~Ug�������)������䉚(�h2Np`-�z��������V�m��
}��O��ߌ��t�M@���ȡ��tˍ��?A�W�7w�MP�j�n(�M�z3��w��e��S�Q�D��$�^�GD�����z���XQ����(Sb�������w;￈��һ}�����w?/|��2fn9�t��m�O�>� |�P4 �.X���7}�M��.M���q��L�f�qM.�|�̙c��`Ќϛ�z�S�@W�mƠ63�UP� �����5�
js4��B�W�x�� _;t%���`ҏ��1/B�ɍvݯ�iM9[S���C�H�w=wS$l����m
0dt���.Z�½�澇���0����ٔC)>Z�m�Nc�v���P#P��qF1�p,�Sͮ��3�g뙓�[Ϥ�cL���'_�5q&�H�(��a��l*�4e_�b����m3�;���2]�
�4�v1G�����F��=����J�1�x�L���i��ilS}� �@�|�D�h�g�?��&Ԥ#�l�vk��|v���(�.��Db"�k7n�`�PH���jt��#E*�f��eoMR+W�se��EX9�a/�C��m���f7�`��QC���%<�Ѡ���kv���=�*���L̝���?䙧�4ֲ�z����3~H����>X΍��Fh�֔�ct�ţ1a!��\<8���D�a�,S:ab{����d���ÒU�T2���������׼���
&F�я˜��E[�#I��Q��[�����������LЅ��]���Ps*D� )d?[�9���ߘ��L���]�nr[|BR�`�*��"�n��?���n��C�秢���!Qk�Z���M&�
����}�ϰ�BD�yM�X�"��av��3dj¡T�
E�V�d}>^ZU�_�@�k+�n�p��N�z��ޱLI׹쪫���2��S�g�S��77̤�ŭWŲ�~v�Ք�f2��0����t]
��a��q\�]��������1x�*�����LN?qnxv�����sɔ�鐪�Dz{���r�~c��-�����\�w���|I�~s�a����Y�?��%3J.{}�l)Bx
%�/��^v�=���ڛūmN��ݔS㱭ͣ�l�٣���|��J���Ħ�e���6��j1N#pUӍNZ�Y��M�5#'3�7���i�᚝�Wh�f�?�-d�m��6�fP7O��0�1�5��Zr�d�H)��[���C!�Q�&�Jp["Չ\ZǟL���>&I�`�
��݌q���K���p���󫗌��ח��mU��\u����¢�y���>\@״QP�>�%ev�M��ӌL�U]�v��S��L^�&SW����M�+�W������nk���1�`�&YNY���>:�Σ7h�JV���~3�\?�y�\*J����ŌWa�bB�Ko~u�z=�_��*tO�.}|�8�eM3l�E=��H�ط�>�U���<����w��8��˰Z'2�ؐ���C� �"�\hdX��*�J���*�U���=̝1��?�?��ϤZ�F5y�\����9v7���\};�);a�R&U͖U�:�p��T���~�Ӓ�� �5��?��d�KT�.U��Z5��]��'WrԜ��4�[Z4��tH�0?���U6-a�p�ǐ]�Z���Y��O�!�"��\�rx#���cikO�s�`S����X�U��$"�s%ꮇ��1%�e���$F���E�Ւ���T=����S�L��[QBUЄ^$
k��#�g^�&�b�'�q�!�0y�4�ټI���;�8n"k�*���Rn}�M�	�|��li�̚:��`��^�e����?d<��� ���z�!�C&[Ǔm!��窳v���c�J���-J�0U/������X7��X��՗O�����^E��qM�%�LNé+Q���9�C9��)�rb�2_��,V,�Oq��
��.�B�hk��l�`0L)hqگ����X�]T�A�T��C��h9�Ԡ��"�����'�6M�b2�����~�}�yw@�0��u�T�9r���/������N�e:3�ökE��%�Ο�����=��7���؅aZ�:iO���?�y�p�w��g;����/H@ 2���3ĥ?9������>�k*��N���]���s�I��#���/�5��#�q��R�F�L
T�����V����M9����Ȅ���M����G���Y>���Vrn���Nr�a����0�5�/.8��i8�{�4g���lR� ��ƅ�<p�Ἲ~tӟ��L"_i�2�,@�g��6��o�Еs�?��r��@�^�j|o���Mr��k%d���LG�Ə�n�hnn����&����ֺ�kU��S
��yL���������x���Do�������x�]��/����C������v=���Okڷ�W>ov��d��j���?��s�}dd؀�F����q�~�q��+���l����任��ߛ�(�R�{�K;tu�z|3dEd>���i��i�.�U���\c��N]#u(��������8Ҡ7����U�yu�s}�t��6\�������7�L6ov�?<�4�b�����T�z)��@%��D�-��UC<
��V-H�d׭e��8G�9���Mf��v�_^΅?��ɓ�Qȏ0y�X�x�!���H���{��^�w�mJ��)�ʩ��F�g�o#�F<�ĮI��P��kM 0�r؃#-�235���?�#��ZdF1Z-��|C*z<�	�&)f3T3���ր�ċC5�J�@L��LA�{���a��&ծk� �dX5<咒��F�VwK�Z��"W�i�U��	75���,iO��)/)_Ѥ���88�6\�R��o���#׷�N{����'xV3�+�;��駞Bט񍐢H�n�#&�$�9��������3(ZaJ��P'�B�Wa���df��"��ÆئXI�6��ao6y�8h�Q\���hu����(JM�S�3�y�7�S��C8a<�5֬�V$�r�u�Կ{	(+��P��!����;�`~xHAE�VGH��ryb�Q8xX�[�������'"o��dI��k*�"����=�{}%���F~�u��-�\��!�"�y���I
��@�
���J���:�4��D(�B�\3aP�+p�����ty��܁j�	a�_��7s&�ɿ}�7���F�M.����Hr6��;���14?��!���մ"���2����ޞ�����of���gXV�ƒD5��]�){���w������W�#O�3��x�XCk������l8������a$�A@"�B�hq�3�;�o�9�r���aV�d(���`���s�s������w|�/���s*#v�߃�<̌h�m�Lb��,]߇=y
#�򛉍�]w��ѵ����$�5%ӡ�MnDCr�U����q��5�+��ώs:FK���>�J��]�22k��E���n]y�ګ�M�n۪�|X^)7T���-�|q]+
�1�/B\낞/9`jz�}'̟�/E���ɾ6@Y�Τ~v�j�K�C�
������;�T�����]��@V]���z#�Ӎ�F��?7���1�;�&QNݹX����ō�`бu_u��4�nrzS��q�.��y҃CC�N�I�SW�}�����\�5e�z�M���Ε˩	�ר]�V:�.fM���s�c�3^��1t=G���i��9�a3j�V"Ѹ��s�Q��|�=� �����A.��&�ۍ7�a���։'}�,�|�B<�2��Bw�����mN�b/{�p�GI��f��r#�&��+~EwN0Ɛ��wο�e<�x�l�Jf�jLKZ[b�o�6h�D������=�JiC�z�K1�p��o����j^�b;�5�[�ץ�1�XS��H����!W�,D������R_�1休l�Q�]Ԥ5/V��k^��E��Zp���&õ�Ē1��M���Tn Bn`�t�!�l��2gl��V+�2tu���>�PV���*n4~��d�H���jI��3;Y�r)�>�81�J%������CH����O�p���J�];&1:M9;Ą��9�X��k�#!�n�/����r���qc1|�0���_�͇�)��᰹I��/7�κ�ŗL���]��7�P�L+���v�0F�&x��{��e���U��8�9rA�xQD$oҥP��Y�­������������o�����g�d�⫹���
D)���x�/���B�8y���a<�8Y[Āo����CXQ��"a�I��s�N9x忔Ļ�P��h�/��9�z���@x�P���]�`��2�����lk����#_��C�*!�!^��C��}���!V��D�N�a\��;��\~�3|�1���I��!�u��s�!{qʡS���<��� �1]��*vmS<z�!n��%\w��v*|�~���XI�V���<��&~x����lR�*��� n4ә~x������vMc�"?	P�T��o��ы&��j��e�a�K��Z#���O�����1р��^���k~V/`��0F��a�7�hqf�F5� %u�´!Ę�f�R�V�H��6dk�	o��6��"���h��T�/0w�[u��$��=iej��D�Ո�n�+�`�J��[����
�(�*3����,����/ ��._��x�=���W/��m����ծ[ݩ����V�⸵����Qu�M�s��4�V�}�@^o(C@'`oơ
����mC���1��M)�lf�7�V��k&�53��X�(O�    IDATG m���W���M�Q�UW-p��tl=g]ȵG׮\ ���o&
�`�~_�Gݷ
�>�a���mz\ӊ�tz>?#C�L�2��5p��/���n
�E{������~��~�5e���^��Y���ٔ�3ad,��L[�N>�!��72.^d��7���}��{�=X��JZ�;y���)�}���?�'��Of��	�::"��A_0J[K����E�+�h��z��8�����RWd�r�uqW��+�����Sp���,j�U�爠�|5���5�.
���E��6HW��K����ı�yg��!�1���%�îʢ�Y����d�����U���H�r��x��!�&T���E���CN��d�@+u��{q9��F�?w�8Љ_
�G�h2ْ0q��rl)�n�@�s��'�3��h=�i�E|\}�UxCaN<�LV��X�m1R�Q��� ��f�h%I�n���7>��gJ�I;�&���*�dI:�__ǣ/�û+{��T�:q�A|ՊёK\/����ߎ�9`��l?!N���)�� O�['�Z�����6����XW�r/�<e?�Eȩ��x����ko����s�l�g����=�n�'ƕŬ�3�|ڗ����qЮ[��3�q�!M�+��Ԫ+�}��c��e�����M�N�ވ$�!���*&Ig�P��-Ǧ���#X9 G��<-��ȬEǆps��~��~.[O��ض�-ʶ�����r}Ͼ��nbi� �J�G�H�)m�pW^}�#>]��`2�p��/��	4���>��FƦ�,�kW6���Q�	G��<�X��J���LfδYL��Uu��lz2����짜R���A�&`���IZ�9i&�ux���H����%�hH���	͑Q�"��K|~qq���9��f��IrE��R��uB���)+�&�V�����4�g�-����;ev�HK�R3�Fx23���G��45�Fmb�����)��Y�:1�(�Jh�D�q�-?�XY�+I�Wk�x���x�-����'�����4_����c���Ww;V�b��U��.]�@U#c h����nV����g����Ԛ�Ju��Ru��.\]pS��3���Ϛ�W,s����:zh3]]�:�f򛎧��r�9�����hԵ��0�B���@����k���:����黦z�������B�O�����Ɗ�H�,�	^��4���y��ޒ��:���>� �g���e�}��/�X�_�H��nܼ^]̽���?;ﰛ�*t�]�q���S���=y���9�Ø0i*?�4S�l˵7�I�8n������q�c	Ћ��jK�1<2��ŎF���ض������~ÈUNv�dP.vU;t�a��YL������A"� ��~���vv��0�E<���g��w��-�+�=��΄1�Y�r�c��6��a^|�)�Lkg�m��7��)�b%	&_�H��3z�X��u�rD⳴�(d2$=Qb�M�w�p7���U|���?���ї~��vl�
��#���T�z�X�(����� 3@̿�-�R(B��3��P4E(�j�5���䴓˦��6�}&���+n$ڒd������,FLֻ^C��K�X�W�Dѥ%)g�%�{�|��-���$��g(`e� Q(A�����+o��49)�	�ZL����3�yf��@W�J~���"L�-U(yjÍ����Ǘ��%���[�D��ͯ�<����J�Vpj�z��
����s��❥_�y�zl�s�^��ư`�Tm;����.3/�B\:��X�	�*g]� �Vp��)[!jv��x�Û�X�#�^v����Nށ����?ZF�C��7�io8Ѩ��*�z��F�AHɗ��)�����a��$U�-�J��1�*�2�d
�Hw_mȼ�C U.@�TƣV2��K�.O}��#�H�X<M�m �
�Lc���9�� .��4&m�}�
n0f�o�-	�`��qڼ	��k�}��\r�"�n|�i�Qn�$k!Y�z�FF���
	+Hnx������z<��,�x�z�B�T5+1�����0j�X���2l �V [{m���.?���g��P�82r�Q3y�ZѩBk�`,qg*"��u��aB��ˏ����PUcՈ�D�(8
~�#92� v A�����P, ْ��z���f�I��'NZ������k��/?x��W��'��"�V3��9�@M`(��:�Q�&XE@��X�+���~MB� ���Gu3�D��Y?kw-�T���\*��il�ۛNo��}3�Ev�u��KW���覉�qJrݯv�:�Σ�7�[>��#�Z������hZ�6���*8��ԕ�SWQ�c�w$��q7�(�<Fט��[[���K8�ϖ�)��=vg���∣����Ɔ��7��6eY��6e��T�zË����-׏S�Rϯg��!���#�aƤ..��B�����ŦM�̞�5��8�"����y���,��pG�hys#y�� �D�b�|v�dK+�7D>�o�Z���E��J�B.�eܬd5m���od��V.8�t���
�b�oy��v��W��j���}�a|�[��CN�Ϸ�B._�'g���������ˑ��g���Ǟ��Ǟx��u>ْ.Zh�`�k٢˛>�Z/�lm1���`_�J[{���D>�#X�v3�}��Q~�����<��9�7�����F����F��U&�V��2dz����%"�B�lS�sb8@$�w�0E�K�e��Y�Ǎ�?W ����$�6��<|�M����α��ٗ��Sp�&*S��V$fX���ǰ�#�	�N{��\�������vN	˧��:u�.�!��аD�䃅:#y��4=7�F"�E����;5ʅAC���P��ÎL�}�=K����p���ɕ!by����W���OOfש�R��K�t�62Ūɩ4E�L����n��k���.OX�D�ZB�%�e�¬/�Ϯ�g?]Oˌ�ؐ��Ɉ/*2f����@�al�V��I8#��Jr�G��g���{^�����'�?�®䱼5B�2n9o�D:ukZ��@'@�T��D�[^j;vcT-s���oN���R$j 	������5D���O�$�L+*���
�l����U�^��nM���5�R�RA2�R�h�U$8��w�mֳ�h7�9���	�JQ.��Q������gg�~����+.�t'�J��J���!Z�m�x��\��288L�il(C�4���V^"��=8"�z=fTȕ	�F�G��F̔+�9��|ָ���K���ղt�e���)x���?q�<���0{����O�?k�?Z�1�V3���d�^�Z|>�L�a�K�����Ф��&����֮������k�{���n�k�TGDI^3�D@%@�&|ɧKM�-5�śIi>��5SִwV���\�q��n��Z��n__ȦN\��ލ=fǪ�]�k�4eb:�:�����s0+KEFsį�F�a�_��kSQ�d[ ��� v���F,|�F�Txhbat园f����9�k���,w�Ä�,^�y\�by��k���۸���X����sv���t�ԓtgJDZF�Ͼ:eI�T{���"��0žO9p��\���0*���ͽ>@,��ԩ�y�W��^nq�/�塗>�J���VULё"�P�TTӀ"��~��v��B)W�
����r���:6AoO�B5?l,Gu�6?;�L��N�z6���/����d����>�^z��Q)-ڇ_��v�yw::��}�_9��Ø0~�]s+��-�������Nb�ʵ<��;�;�3�Fqm�j����L˘N�V��ծі�O���WS/	�����:�}=�Fj)V��	��8�!�Ck(�~���מ�p[̙���&֭���h4�ՂC5;L,�����GK�;\~�uxb&�ܚ�#J� D"̘��쎤��|����W�b�jv̞���{�_vef�iX�nI�<��u���kV��)��($rY�J�j��U�HP��ᘑ�ie."����!)�B��X��8�-�Ҫ�MXU��[��ϼO�e4�x�lU��>¾���Y�_�%��Q;�6�~�8b:Vo0@8 ���V˞ ��O��ܥ�e�\��o���*)G�
5�N�`<lv�W��-�j��8��z��4t+�n�1����2|��I�)��Yc���}x������<N��g�����mir���Oi�\(��7�C*B[�Q*�������O$�5��67��R��+r��"52,/�PЌ�����4-�E�CFn%b��2��BG��R	���<��6��%�29�䧲�S*0yL�\���>u��?��D���xjy
��d�$۳�ӿw�8pW<v7�̝N6_4�@�'�,{^|�z6�q�~���g�xK�X��k=�D;#�I��ABn�y���߾�P��x{�R^{�e��OfM��#�x���7r�i���=���w𷍦R-�Ե���>*��6�zƤ�[��B��p�Nje��(��
�5x��9��[�O�n<N�ۃ��6�h��x~e���V�j��fz(���Ó?8�k���Q�=�%/ܻ��?�<�JQ��k��7����v؁'�z�����&�Jj�쀛�q3�\zs/�����E"�i�m�&}��F���r��խk�-�ZS�����&+]]�:bu��қ;w=w	��6=���<�6�7��|uN
~ z>����ٵk����T�x�Ű5�6��iS�ፈ]?8�1��?Y�?����uz�n���ƻ�{��b>}���W�N���`�L9_������s�6ʥ���v���g��:��sT�6t��p��,Yއ/5�W?X�K� 8��H�oHk��C,�B<�P)�͍0v�$�G��e|��q�r�E,���C��[ ��g���@�g���@)�1ћ2��3z���{�S�k���x�~ҩ�f�X,f�7��5x��f����_X1��t���k��^�]sX3\7�2+�&��=ar+���N[���_a|,4@֥D����_��IcY�c�s/��o�������fCO�ѡ���$*}�y��8���^���I]�3Y�j��߾����l�L�6Ր�^�=v�� ^y�ƌ�b��s���Gy��8�S):uڔM�Td��M(��)9�H��{X&�=��Q��yI�!U�����1{O�=r��9e����7S�{L����\9pY��ԫ�����9��{�Q��>�?���zo)�q����D�
�����1ݑ�v[�"0����5�o8���@��`��J��*�Rq�W�X^?�O�f1�E|�V��Z(��D�Z �gu~��xm�nl,��U�첅��J˯���������KƘH�6����#��L.={�Bw�I׳Ŗ�X�;���%�
�(v�g�!�K�R�V��k�`f�Qc:��I-�	
3�)�H&������X�C�##x5�R^}Y�!��Q]��y<F�EL�[*Jw�+]A�=M^� >����8�k?��o���s�C2}�m�x�z^}�=B�8Ձ~�G��Ǉѷf)��y���.V.�-�b�n��ѻ2}�\�N�X�hzF�
�����d��l���D0�a��q�/�OW�݃v��'��Y�+�����ęG�V�F���ݼ��ۜ}�|��{�bh�����	�	�yi^K*��Q|C�u�ö�k�*�K�m��+v����q]o�u�Vz�IF/��wv���K�,^��1]'x��m3�㙥k�}i����>	V�̏�#�������u���C���׶�;'IEl�_�&	Mo`u�"<�ԕ6���K���u�dm�N����]ݲ@_{k]���
���frZ"3ݲ�jW�m�w��W���!�l���g��2�7k��oZ���xh"bѫ����<��Y�v�]{w}o��^�]��N��o�zU1�Ŋ�x,?�h�B>�S���L�3k��5���������H�����~�-Yøٻ�6���7�p��Z��\��]@�N��'���.g`�{�/��n1��p�b��	<��dsun��FO�O�u
��D���H�JF!)Ba?���-�T�(�;/�d$3�]�r�E^�cg��x��L�
��T�Du!����aʖ��O�"Z��Ts$S�e�Vk��y�r�Jӹ�IMQ�>�����!�S�Xݓb����I���%�c�D�e;_�-�pЂ-�ez������Ͽ�1O���-�����ZHn����Q�t�k\q��tvN��Y�=7�IG�F4P��0���'v�}W�L��h��Ss�T�Ɩ2�Nѽ��w�^�QG~��T�`�?���Ko}���T*u�1ơX��V�k���(�-��5L(U0B'�J8-g��Y��]h�hp�2���\Ȥ�F+��5��a[8�F!���X�T� "�1����	���^�s|��l'�$+=�$vQ�TV��6N�"c��ʎ��.3�r�����̘)�j�"-^���~�Ix�Ғש���^3U(��"~y�K�gQ��#o�폽��MU��X*�$�l�h2e�j�%��k �ǀ�K��o 0cx*ZR1|ղ�z?d�mq�7��,N>fk~��%�l5�?��[���H��{�%-����ʡ�8���z�\���k��VI�-�]w���y�hkk5)��o��Q�<��s�1|�b�|�!Gq$˗��{��_�7���2�T���ކ�����1y�$��������3���el�͎�2U�֮⒟.��G�e��l3/�.����Ǜj%�HS��)���on;�ߝ{�)b����>>x�%��e�]���;2k�ԝ(y�JZ�|����|�~�����#�l7���J�s���|�)W��X�ܮ�_���!�^���x��ט�b�]�'������Y[�l��qW?��k+�Z�h�z�i����5�$��p�m�[9���{�����-��pʏ/��?���v͍S_{퉛�;|�������/������ix�:�.?�����<���c�+o�Z*�z�n���͙���}4�>ް,Ui
0�ތ��+U�ݪkV�l�`^�%-в��h] ����Z��^@شkm��T�
��xi��:� Yݶ:a=V���4n�����թk��L�̸\ň��4�Qw�μIh����z�:���t�[���i �E���A�q��k2��s�k�C��2�}�6�2Q��\u+�ѣ�9��0~�9m����7�*�䩜7��!�Ht����%C&�*��P��sv^����{WW����m�m����y���g�}͎n������3x���y����H3z�I��'[��d4�K0d�c�O�,\u�9�����<l�Ȩ��F�MLH7j?y��c��wO��c@�bI����*>+J0��fаo�C�
��b�(�e����	*�ԩ+\7��OVQ�ϚKd\'���q[�D۠\�ʮ礃�������_pѯo�e�B֭ZʝW�������,�\�{���M4#��'n8��*C��O<p���j�#3�5�ݭ�$������?�����}�{��
��Q��r�/�#2e7֫��
}�)���F�����RF�w!����S�
6
"�����"!�7��	�Ì��8|���\&�1Ѻb��LO���$�n�H�!(� ]P�>�>���Y��/O�����/�H��6;x�֘�T+��dhI'(T�T=><� u;�_�*�0��[��\��m:�tA��f�d4�bB{�w���~/6_�c��fϮ?���푧xou/+M%��"'3Ŷj_�^As�W�~��3�r�lP���NIg�!rC���1�J��ky�:��چ�n��ܟf��nz��`C̻������{S���7?�yg��S/�'_,r�3x��a��F8|�I\y�s���E��ֻ�g�ݶcF\�����#���
_|�%G��z���٧��_��wܞ������6���9��?���OcІg�^��oi
������y�ŵ<��+tLޒ�A(9ʬ�Z�)zzh������\x�^�$��+�˛�=����N�������i[Ow���Oh��ʫ�s��}��3��������Ȃ�^[�o���.�1sg�8���������>��t    IDAT"�&t��ܙd�G�����uyN�ݣ�L9R*�X�z�ƕ�͗0J܌Q9����gz����}۵7��\�=d�;?v�#��}��O6�m�8	$�\|Ğ;����z������ ���#�����H�����[�dI��%p�}���]ի����U�g�H�!C����a�u}�����������7�˘�4��J=cҲy�/�W��Y ��R�X?�l1S Mt�_����������Ir�CE�Fn:�
�]��&�N�x�w��
��5�o�Ѿ�oz7�:��Qiy�W�fe������\|��s�	����ˮ��	Q�v�ن��x#q,���U��/��x�U��u�k��N|��0g�LN;�T���5��7p�7���5$�O�g����ُ�v�H���ps���$d`�p+N��%�(d\�E�j_+����T�k�v�fNN����
�lD�C�P�����	i)Ñ�ǰ���e�D~i[=5*�\#��7�0ʥ�@ �Z'�L�%��ż=�c�]��GX60�������#*k��Z�<x6�~k>+��8���	t�@�8��;�E�u�tU�3y3�:m��Q�����@̭�D�*�̃��ͼ9лa�@���?��sl�l���<Ɖ���4����d ���ZcȄc"8+Aأ��>j%{؏?�0&>2���J�e1�������%��F8죦0�ZO~�GE���r�޻����fת&U�H�=nl�\��am��s�~�3�/am�˰'B��KI��HdY6���؛�2�*��/^����x�$Zp39���2�+�>�Oa�9Shi�L���r���!�ifP�C�$w�����X�u����ۍo�̈D�tEH�e��Ӕ�ES���6Z��5�#�����ăJ�y��T��z	��O:�����-g0u�h^z�I���!f��G��oϺ���֛�x����Y��K�y̱�㩧�}��᏷�j:��S's�=����_����N8��k���Gs�G����ظ��Cݗ<�0��[�i����3o��3��;ﺃo|�`�O<��~�z�y���56MA|�r�5�I���_�N�Xq�L��۳#l��Ũ����S+ob�>{���i�ib��!��u�;l7s+>|w	�[��@~Е <�8�/���/���?������ңy��י1��q]����kq�~���鏇�����i��SS�F�^5�5�R=>�R�Pv���Ӗ_qǼv���λ���'��c'��������̧諶0�S��#��a������1�O=�������x�.�pJi����ZW,`��J#w�@[]�@O@'��@��x��u7G����f�xÙ�Q44�o�R���@����~3bW7����s�A�	�
��+���0�)oX���9�:Th��Y�$k*T��8�*$$�{���$@�k��4�ҵK�ް�maCO7�Rٌ	�l9�U�V2<<b��T��=�6q2���紌�����\v�m�ɸء��˒���Q,�M ����(e��}��U�I�8j�i|���t�����_��/ϸIS������ �>� �
�z���z�k��,Ѯ��۴�Tf��H<ָ�����&�>`�������T��(�����Ł�v�?�HD���h�P��$�q�%�ՉF��S�x~�B�%�ٯJޣ����1��u�ft0	mu�����DG���K!��obm��7�6y��B~��M�h��q�����F~x��R�Y��\u�.��`��6n~hW?�*�t�d~�]w��ʃ�ȏ���z�ｐP4Ɔ�Ac�#-z�W��7���=��q����s�9�(��ó�y��>.�ݽ�:氩R�"Ɏ�%MS�g�*xJ�d� 
�R62:E"�Q���P8�#�[�OE�R `�FB谧J-7Hȩ�{|t:ńαTKEF��Hv�r��p���e�8ވ	k�Ǔ���'�#5�an��+9o LM�S6�r�$�\�n��T]B���z/�3��T	zʹ~����o	G�1i���Qm�vY��c$w_������닀�� n(A���U��2n(DM!����o��5��e�"�fg3��mV;7^Fs٭5��m��u�
���W���n�V7��Mh���;]�+���p��HG/�Կ����<�y�-F�W�+�WR� eE�z��1�5�c,�����p��pd�{_�5�[��v@<�zq���x+
�'���g�K���wL�o�H�uz�J���$ੳ���d
%�6�W������W:捗�d����eICO)���>�'+{8|��8��yWd��\y��8����h�����!�<������Z�Ӯ��։ˎ1��e�*������Y�݇��ɏn��5��wA����u��=��q�^0�%^�p3QN;t��wl��������&@�~�������*��O�PP�K��Ԑ�/��7��PC�����o�u��z3ZT�)�U����ak���@���U����6���yH.��U{q���ձk�����i3��6���~�:�����yh���@������n]�oj�5���4I�s��й4��c������W��I�rF�j�����m��}�F�|�W��Ц^~��K���U"��wM>�����	��Ʈ5?���X�^���1�%˒w�e|{��t*[�۞G��'��]���z��M��<���v��䙷���ڈ�ia0�1�l�w,�C$jv�b���	�|O{�6���J��`(�SظҸ�͘6���ê�T�$S��CRf#���5l"��.���6�#�+4���+�0.o�wX��P<h|�i��:�ݫm��+֓�[�L�+=����DH��qG��]�NZ����o���3��KOd�?9���p�/̺�ǿy�����Q�"�]u.��B��+������mq���2}�,�>����&O�"=�����N<�lz�yF�6mc���3������T=J�sq\����_�tz�9n�J|:2�'��-;�d�T�ױB~*2T1��������Z�l֪Ec���4W09�UI��N�3 j{�,]��>i �������ު|��~ꎒ�lc�5a'!J�׬,�v��0��y��p&�80S)���Tר��Ē	�#M�'�c��W
&�Ȭ>�!�њB�y�-��G(�rD�����xO�F���\��p-�l&�5n������g�O��5����U�� u��M!������B+��7%�W��E���>jx�a����qT���2^��*u!���x�~Ő��� ��}��8���QðI~�����D��W��}�qJO���QRK�{�H�o�#9��{-��(�z���-5��9�W_~���l��3_������=����ͷ�ُ9�;���7?���SN�ct��v?��'r�;�d�&����Q�"D����R���)ej�NU�5��������sѧ�; z�ߺ���8y�s<w?���1��[��m�����9��ߏ�� }0�ʃ�en��F:'�dp�h K %��\]��ƥB� \s.��M��j���Igz����A�f�Zs�ۚ&.+W�0`�Y��N��0$��[�+�U,@V���1�q�BA����������5-��K�C��s��M�VG�ק��h�t@�RѢ��z�*:���v�$[��г�T<fG�(Wl�b6���K/��Q�&��/�Y^A�����=y�k���:&!+R`Q�y���
?�6�)��F&�n���ʤi��J`�n�{o&I}~���v�ݙݙ�e�lq� � �	n	N� !x4@����6��Үe��yk��{��>���\��~�}f�������s^9�9���7ޅ����QW��͂㯅���^�,�d�TWBGbP��#��Mz�<L�B>��v+=5?��v�s����_�O�Q�����p�>аmO��s��������:Vs��F$X�9��M�X�'.�T���s<ڊL1���l����I/�#9��V-�x3*�8F�{1kB�7���|�j�j[.�C=�x�����0y���ːHf	��s�M�L���Ȍ�!�a��r\��46�9�S��\l��c��ŧ߬¼-w��.B�T��;�`EoJUh4BQ�q�%q��-&��bj�z�U4vt�q���h%��}p�1���Y6DQ�-T�b}�S
U�8� D����[)���PjeZB8�\O�9>?r�%�eW�R����񺅊�-�ޫ�ܧ�r�5A��s˂R�C���I�ï;�_�(Y�P�^.��/G�\@@��G�,ǂ�TP$�.AآaOnL��W�Rl�gei�⁰��(�I�s�s3x]Q	�B-4�	���%������V�%x�I@�3FO���rV�x�<��'*�#��|��$�d�>nZ]��B���z?������j���Q٬P�V΁���7�1$p(Q�MW�U*ޤ��_<8
�k�u�*�����n��c9�CK<��
��#��2u��#�����F18����H%�2�>�ɢ�c�ȯ~�n("�"�8�k����Oa*� �R�"�`5�#>YG��z]�l���RC~՛�*�u,��ƅ7?���s������b Wx{�>���}��p��8�}W��S�����>��� =S��S����{��5䊎 'A�:g�Ҹ��4��BWU�����u?��̜	rU@%��L��ٟ&����B 0Vi�DEG�@%�VMW2�3n���	�b>�|����RƯ,�s�#�W[ �Ыs�U��^����d{���Tg�)�S�����h�Z�O��D�hnnD*�D����H�Q[CWg'.��2�wNBr4�s.�-�n_#>Yޏ�R��	)�����*�������C����@�r8:��k~�t.+�����5W\}>_�
�~��Mb�Pe���E�!�Ed�9T��7fbx:��"J$e�U�A)f�\sx-�9dO̝֊瞸V!#��B��ü�����E}�����E-[\T�N�NL�>]�?Ɋ�tF�=y��Φ�k�f5m!~�)(�[q���`��ڦnX� l-��?5�9ČӲ
��څib�w@綉M(9	��YT�z��(�c��%8�1� ���?��j74t�u 3�@�@�0�-�X�7$Y�j@���h%�(�:�p�[l"�"FB�q�����(�/�﮺S�,�^����$���H3J~S�8\ݒcW5��BY����N*���`��B�-I���-(��y�n:@}��d�%�����*:SE0�6�L&ݤ��.����b`��R݂�?mjz�2�Ӂ��5���:�]W�s4�"�P�J�^�@�j{��T�$�5��ꢊc"��ܵ�T���\i(���xM�~�-��6G�DK�v	�,��
B�q�����Գ+TrcI����U!�pꄣU�쬖Խ@�+�����^5Kf���:9���9c	�K�M�� E"cՕ�ku���p�� �ߪ���+�;J����7�hj@Q
)46�*�FG�ŏ:�1
��(�0�L��G#Ru�8��V���E%+wTh}�jO4 �ЄI?�b��/C�D,'` W�E��n�a�U��P�bٳ�%٢乨4G�m�U���L~�{.����4��񒥻q������Q�����U��>��}���D��'K��-��߲ɹ|��b$АT��:^���g���$��8�����?�~���8%���%�%HwuO�' s᯲�	�\������=�����9�ul4!7c�UH�4���ZZ�xd�WU�(̢�7nG��g�*��=x||����s��^�X����QL�&#)K�YM� �N�{�3Y�/��ֆ�\�D���;���x��%���P6�Л��� �s�XP��=bj$���ڀ�t��=fK���֊�?o��:&v";��v�n�{��bQF�-Ob�î��q�(Q���h�'�s6��:�4G@�<�dQ侌�5~�Z{PY���
hv��t"�#���\��>?�{�DB9��쳏���b��r}T�-m<�mڥ������ �=�q�PmL���&Xe�,��A�؀��k�������vҼm�_E��"!� �.B1]��4F����;g!��a�P|��P`M�Ģ(H����AU�7W:Xy�8y����Chi�Mw���j��c�R\��
|ao��*��14V���NMp����k�Ì���1�%���rNx\]G������"|��-�@0ڌ�F�U	�03��k�� ��+<Q��P�8�Jb!'/�od��eOi��8��8R���L
È�e7`+A8$��ӨW�G��Pq��=+~�80(��A%�CQ(�F�4k,2��p�r���QA$߃�m#��'�+'�3D6����jQ����5��:�cfNp6�mf�4�d)܀K�5��d Ev u<��2����^Ϝ��vø��Wq�I�L��qES����o�Ⱦ���j*B:
C��I��*�op���]EH�l��H����
:�"���א�� V@�h��}(�� � 3�G�GM�	�t�UF)�M-��'\�R� UBNBP.���c̲Q�l$'�
2%
�x�^����+�\=5��W!��s�[��N����^��Z2� ]1`�a[�mVSG���]~�������w�;xϭ���S,O8�П=�gH;�������Г5�=�D�%w2*5Ǚ��z���/JϹ�~	E�@F�#��A���oK��ź����6�\��$�����������eyf�[�~�\u������1����p{����ex]3dF�:�m��jY�`��s;'���k���c��ٯ'��Qe�30 ��Ҹ�9}]S���%�`96ښeX�����2M̛3�^���a�����X�>	���H>_�6qS��Ξ��:������f`�M'�³��}��k{z��Ԃ����מ��+)�I�K7�qĩ�"�2Kf�)8�tDB4Y�P�/�6|���c��'S@���w'	7ۋ+�;}��o��lrL���}�]зv-fm4M�����P�o����H��N��|���EOz״��Ԋ�i���E���� ,�Ǝ��3.�O�ދ3/��7#��!:َ�C�(;y�5!��X9���Q�R�
�,P�V~G�2e����*�����"�� Y��ԆD��j��`( eU�>��?�����ɳ_� -&h�� �T��iQ��Ql3]Cw]���9L�<[�ޥ��p��vEE(L3��0��b-�Y��.~Kr�h�Gg��/p%I ?B.��a/~��|[l�Q�<ys�F�\1�׏�����_Ǌ�"�m'�=�۪FX����%|�|;o�%~s�T���]��^yw]v
f5���>�{S�&��pv�~\x�l9����^{7�H#N;���k&0P ~v�K����O�m5��+^���[|�vf�i�٩	5�Bpm���=@g����������|��0k���q�n*�:>P%��r.`�q><e���}\���VV	H���)ñA�zS@5xl��ىJ!�;�|=k+t"뽇��pb�^*`��&7��k�drX�d-rY�P#ң�}�9���l���`\��J@C�@�C�~�=�
�h-2�HN�1��SE�kod�)�Е0�no
f	n�/<
+��?��r�܊���\Vgtj�P-�eb�)~�*�v�M\�=��?�����M��n��^��Q�tı���W���������/_{q��8:gS��cfX$��ؠ��0��"��쩲���M��a5��L�:A��kY�gVβz�&&@P�N�>�|uK�<.
̖�_����0p*�UP����jɝ�WG�)V{�����|�$�à���f�UC���o4K��Dcsڛ��j�
��>q1��Ǡ�vu	��O���P
�\~3V��a�ZГ����1��o��U���)GV�/Z    IDAT�^M����F�&���?��Ȁ�x=���	�i�-�t�z�z��X�o���D�6�XG�%�b.jk��+!�G�R����V1�lbZ9��S��K�S���_b�'�@��0��nI }���}��K�D�l���3g�w�Ì���kٰ��s6g����~���b��9�3fnE���w?@>����8���q��O��G%����|(�I���l���J�~h� 
�l���yv�hFm��RJ�}Vυ�/����hM�_�CF��@r�.qf�����|9��d��暺�R��t��|�����bc�M�cj}#9|��V8\j���M��"׿�8pG���LO�O~�[_Y�Ps;��*\z��8x.��]�2��q5���/l\z�8tׅ8��]%i�x!����c.�Fi\t�!�q3
� ?��~|���m,�N�'/�����w��C���6�{�}9�Ș���*����c������"�K�c.�����\~���c#�?����ݏ��x�׻�<�[�~J�z���u.��Q�[1�B7�u��
bq\̸=�&/���0�����-�s��WU!�}�~�oFpe&.�x�y������[ao�ے�w���c ?�:�˹����8��9(����3QD��$�Y�;�J�\ȓh�(0��;�2�2�F���7�F7`��U�2k6F�,Y���Wc�sq��gï�X��Gx����8	)N#-��}>᠆{��W����@�G�°��i����`U�6���C3��P��I�j%/V�����:ku�#�9<�� �y`���\p���_�}��O=�l�v[�{�3/�5Zq��<�]H9��������S�_��R��+/����E��ʪM��Uk �p���깗<cfr,���{C�BQLJd�DS���x�TZz2�`H�Ez��`�<|��R�����DJ���!y^T#�1��z
p�R�۬��N g����Y����Ep{f<~1��x^��l*+����]�Z����OV*���}@0��Yn'�757bph�PD =5:ۦv��f�R��!%�=�Ԋ��$ξ�wX5RF�hAN��/càa�8JYP��E8��\�!��$�>����� ��
�'}VqG�JQ��@���.�%�0�;dc�Z�$��9D��Q�K�"L��PX�_� �����o��3[�%`g��¹0F�EY�l��n;}����=�kE�K{EZ���z"��߫g��Ú�+Eݬ��>_z�l@GS����S�z��!�	N�dX�z��Bi@��F���2(g���0�=��1�ϝ5�D�/����Ua�
�O��m7��D�� YN�L| �[Q��ա���b9(d��ku5,�b%/�*��v�]F�F�8�g��}��t�A�+Z0�02&K��p��^A�W�2���4��N#���r8�����ճ��ѻ�9-Н2���%C1��Bk#S�#O���q��G
P���2|����z��a�F��*�.��'��w�#`zܥ��D�v��3����K�}�ml��<��L������Qx��%x��(����+����ĥ -@ҿ̈́9V��>�����'��k}vٸC�"<�v�z��8t���>��'���Oq�1?�Ďf�;醧�����V[BA�����9Z�1����DF�x�^7�uܥ��a���K�inW}rЅ������2����w{�6�dܜ`����+����y~6�|����ȗ��[�p�������pgQ5��Mڣ8v�V<y�������c�8w6�YLFq�������p�\q5��c��1]FZ7�~S�p��H��&��|~�3�N���,�O��)����Ŋ�|	��9�f֓��!D?��Ԋ�֥��޿M�}���e�E�o��j*�\~�ݗ���0���^�r�W��]�<�7Ԅ�p�a_�c\��?������Ñx8��_��I�H�3aq���,�3���f(��� ?<�� .=�̘���ڂ��F���� 	<�bd�RV���Aػ�z�c���[���3�ol���XN��5��CKk	h��d���0���DG� �����Ys��#� ,���I�"
ò<���D(Œe�1w�|�2Tg�Dq\Z��4�4	(��]�/�N�������sVڛ�P��i|���:�%�}<�U�^���6�H��n����P�L�)b4����[�\�9ą��#�#.X�f��MAwM8�)%콖JE1��aT?|F�A&�=���d�e��À!}yݰ�{m��`^�.Mw��=N�p+5�4�_�~�c�p�o���d�6���.,�77�bѢϠ���%b�C����%+���G��i��p�����5ذ��1!RZsߟ�ՙ
.��~|9\D�u�̆������zDWF��bV�2	Jr;��7ˏE�����X$5����/`�����ݝ�nۅ�ooA����*����d}]8�2�-]���Vª����_Ǧ�m��)3�����}ݢ��fQ�v@&�l�=M���0(S�ܪ���8���uM��%�{�8	m>`h�(�:���T�޿��L�?�&W��4EG��a�>g@�Gq�yGa��瀊'�u�u���_xU��{�=��O��]��zV����C��qG����T����79��d.n;j>�����O_����\�����3x๏q�ï!�1j9������х�U�K2^��և��FS�ߞ[`,v�x���� zS�Wޏ��a��<�v��H�����;=�r�͖�6��AωХ���ϗ����5�&�%2��t�lɆɷ�x>��F���i*x?�1���׌=�������H�ǵ��Q>��D�.%F��`2�9��4Q`�M��.f/�7�a�Z�=�EE��tM��YęU�=���G�����v�u�X��bl9k&.8u?��L�Ѐ_�z
>y�E�f�����E��B��޿o���<���n�d�P,J0k�G�c�M�|��π���l��9n��:m�9H��N�E�g+��T��A�1���Q���N��O��W��!]���+��HO��q�O��~�������{��+��+��}������V����T	`,+SUu���/�[��9����o�z�ɬ���̄����Ԫ
tU�4���\Zcf�	ScPP�Є�n����#=�'}�t>#G0^��x�֬�On#,�|QnX���ӧM���X�l�K�	�Ϙ�b���фl���,�r29�p$�h<���A��5:"��[�g*���1�Y��,�l�����ճv=&�M�a."�HT%���GȇuX�����N����M�pN�Pʳ[,ҋ�'a�
�V�nW�7|R���C��Qb�N�k������K,dХSW�K�G�!�Hm���BҒY���+�2j�(dJbDA�u��T�U���#�j^'�D�Z���?,l~Jw�}g����)�W�q�Ka�ͷ�s/����)"-*��f���g�a D���Z$S��w�\v�Nj�+��8m�M�[9��	%_j�a�h	+8������(���3g�'��[�����Z��+��a���Y�~�kX����\w�1�[�
̑�l��f�S&#o��ПĎ�l�s���hnh�c����K1u�B�~σ�6gcl��~8��{��:y���:�uh�Q1c�,������;,�F�OOs�Hm�A!�Jl�>������&���	'��0(Q?�!^^�T���<tO�8��3�8릧��5'0��n�)����mQ�pщ"#��KKq����מ�5�5H�����'�=v�D�����{yl��<���-�8|�}������k�5���h#���M�D���W��'?��8��j��<��9(�([h�P���Q!�n��fX�_��_�;n��`頍��|��q���q�1;H�����'ց2�5�H��a��-���^/��GH�>�ǳ�*���>W�ɪ� ���d���=|'i��yΝ�	p��"*>8eC*9j��|�Fď e��kT�GN|�`i�T�<2���^�^ua8yq��TL~�rZ&�V����=����6�nd����E�XD�,��$��FsC-v�v{����W_���4���rD:7�>[��ڊ��#�^�||QMK")��ӉG�@�P�pK*j�KZ+.��'$3����e�QLK���6o�1%�����~�?ϗ_~�|k׍�܏���M�C8��]�+R��/��� ]���?��r�-�x]�x��-�e��d�q>FGǼ13���|r�W%Ty�03�0�]�gIz���"[5m!�13&���_e�S�%�/��I�^��(��J�d�h��Dks=��fϚ�e+W"ZӀP��sg�$�E0���2���]"H1����T�*�QW44�����r�\F<�Ñ��}GF��o�4�7����ud_��^֞N�D]�>Aפ���h
]]ӱrg��D��҈˯���&�ᬋ�Go�A�}��֌d`�!TJ%>T��$�Y�2���5��)�X�{�EQ,��ED�aME>T�=<�m���vj(���L'5Sc
&�_CM���D���U*@w*����Q��#5�
�ΚP��²Ma�o��Bd3#���"�X,��fm,�O=��\O��P-]�L�u����db��j��.D�5X۳A�=euu��cĮ���n*LLش���:#��~w
�5/��!��{!V���y�o�G;��SU0�^Z���{KLWB��x���0�͕�����z�m���.�w|�j	����p��������b�Z|�/D)�X�P��������6:�ب-��� ^�˫�>{>|k�d$�Q�y' �<[P0(����q��Ux����դ�V��m7݀3�8���;�s�ojŅ'�}��qM����A����������݆�v��+O;Hz���c��ůQ�Ǖ���'5"i'���>�g�M��v��w��Lӻ;��;K���{?�+�7��ЎԆ8y�i8��-�z��_|W<�"�a'���&Sp���
��K8�P0Q.�7b�P'�{y�7��j�N���S���Z�q��(k��}�?��I�z(�L>+�*�-��M�x���!�\�����w��}�9нҷ˞���U�pE
F^ʹz!�}�l��c,�O��Z���
6��.�䉜�7��� S�m������B��d���s'S*��o��
+e>�r��Roa�Z47u`�`�X��A$3�@q��?�[L���tj�h�vu�O?��o-�S//��8�H��Ӂ�ZdJ.*�O��������E����檲�Zv�Kb �q:# E��E�^A:�9*�%~'~�(��:pTz�Q�Xت���^t���]���	�.Y��u�p����XZ�k�l=�W~���������P�RQ?y��o�����<c��X�;�����_I���n�a�UB�c_�?9�����Tu�bFb�)��Y'�-m�Rj���Lgl4��Hȭ5��VѬ@�1ir�H%~�����B��B�yD�PB[K+r�Q$Y�
��>A��ں:�R�}ڔ�X�a�X|r\kddL��hP>++�HX�VS���+�\�%5���*"`�Ng�vm���p8��h�T�I\��2��L�L6'ĸh<�iS'㪫����Ã)�rίQ��#6a6��fП51��#�éhP]Mz��+�bsFEѵa���CN</)a��3¸nhj9�|��x��TNƄ�j Z�@$��dk>��V	@7j�\�YR�g��.��L�*u	(�a�y�X���x��GQ�
3�cJ����\B }���4J�����ko`�9s�Y���c��O� ���ï�\���m�@8���Q�"�.]�ϏI�fⶻ����dp�WAk�S#��U�p�ŧ�+Xg��]}%&N��Ӯ{}�!��<l<%�U��|�M��6��_�އn8��t\��A����Hw���1�57��!ǲ�ze��hb+W�Þ���7�!dUw��
�=�b��b���6M(���k��7����o�7W���BY��yj�W�W��|�bs�����0oB:��,ACEƆ�����#e�p�9'c�i�2֎���C��Q�v|��bA=�?~_�0���qˣo�{z7n��`D5H��'�_�_�~4~��LY�N��z|�.�]w�ם��<w�]�᭯{Qd֖�ǉ�o�s��M ���_��O}�n�0�O��n8g����8�����c��v�P�����X^�Q�^���-
�;V�	W�I���?��b�z�ß�޿/���S ��1�� ≯������:'ĭf<�����L:�n�2�'5�v��O�5�9K��$xVx{i�0�t�*�-�bڤ�=)m}�����:;u���Ě��1c���c5���4�i���KR8�i�P�����
]˘�G ��/1�<G*K�����L�����	���[���ޛa���'��P&�tH@�|�W8��S�j��W��ُ�cU�Fۜ�K�`�<G�`LG��r�_�}Ώ�����E���B ~V'J�l��U�%��G����Й�)���cn�����殹�S>����?���/zs^�f �"�P(�ض�R��I����/��� ��������@�c����y�Psfߙ��"��w�_Ha�P	�̂���e�c�&�I���Na=k֊y�̍�cpd+�-����V���DRԇ�������2b�Z!��%Rb[�RG�@�D����`}� &wv�*�D c,�BCc�$���e���+������2n�W]�l��X�L/3�c#H��a��n����k������1w�|�}C_���Z$(S7�=�k�btxM��Dhn��o��12��)\�Y�@+�f��g�I�fO9�M�pR���ȏm���6qLIX��NC$�*������>tMi�ΦV<���0"૛��b	j��X܏
gS���tѥ�!����JT��J~(a��m�r�p�I�ﮋr9���(�͝� �IDf%Ǉ��֠��}���V��Hn3tΡ�%��3�)H��5ԠP."�IR#P��S6G)0ϼ�P;6I:~na ]�n��Tl1ч�H5M�x��\~�k�Y���$l�q/Ź7܍D-���ќ\z�.�(eE���Į{쎥�V��T��6�O�WO=�4��|!����6`˽��B!d��W���^��y���d���.��7����^�z9�dC("
��"2��/ ���;��e��@��Dg�F��
C������_[�+/9�L�h�G�y9.����"�Or�/�����h�Y8︃�H�[����`��a��FQ{��,n��.w�8���`����,���w����w�Snx.Y��9�z[vO���'sP�W�ƛ_�BA��SϽ���g�tca��|��<���:E������C~~-���Jl����x�S�Z׃���!�*�I�=�or~$�(�B`�͵�y
���z���+��[�=Q���̿����w�g)#^�2�恬��TO�U���ngl@ښ�s4��GW���/�K��o��&�>�p�m�y�S�(d��#�r�*������q֜,}Gc`�`��?4��3�,M���!Ģt+"�����P1�#���/��U���b<p�C�0	˗|���xw�u�P��p�q���j���K�w����V�������|4	b�B����8[��\;n��A#%�R��!����]�����z������N��Ǟ���O{��W�\��g�;ߌٳ�[k����7w �2*�ԛg�P��������� �x����z���nE��$����ߚ����$ٌ�QK�CC�:e���i5�l���蓠ɑ7��Ŝ?ًfO��1��<�
zĢ��S���(�I��O�^4IoS7�E�Ԣ��ڸ3@. hkm}�\`�%=g3���/��δD�    IDAT���R��������丆�E�����(�L�I��V������9?j��3I̜2v����~q_c�0�7���-�����}m�M����F��7�,�e�>��L��\$�5\�Z&���}#|�� �E5�8*Nc�^L�֎�=k�`ތ�x�ѿ`,k�_�V�Ԡ䏢���b�BZ.cJ���v*�s%��6Xr�'P������z�,1g	qD�,!VŦ6ƒ/?G{k�G�t]��Rw>��cq�"��D��W_I��j��r��ｏ��z���7����J���hh�%Ђ�� �r~�5�L�e��W��㪳OĬz?2#��j�������@����P�;�#���y���2��03^�o�9S[}���l����o�>?�_�bҙ��ls�7�㕧^��9s�ʤ��w�z��J�խ'����w<�J��W���
:c|��稭mC�����@���ۘ}r�:�z;�+O��oṚ�~�3X��{m5���_,-��s��-�\���xd�{���������}>�9.=��qtH��7/�2z_	8�̇1��c�M'�sw����S�x�{��/}�������x*��?J�$7��o.�{y=� ��$9�snyo��6��Ll6#"����cϺ�����FX󎉳�,<s�׿rq����Xۉl	�7v��̍��Pɯ$�@o� '�3n�V������͏g��+�w���.�b��-�2�.�@���e�^�,h6�l���H��<T%��.8`'���=x��p�9�S���/�`C�6���G1 f��fI_���,��#o��\�𹪔�Kyާ�iIA	�zG�f!�wd��рCw�Zy�L��﮿_/�]���BGk�<�l��]�M��<�*^�x%*�0�u(�mDkj��[SD��M�j���h���
"[m&=� 'kd�_נi�n^ڵG����0��T5� ���I�\�2����&�0mRӫ��;/�{|�re�u���jY2�f��a��P-�� ���yN1��y����/��� =��}�˽���Z"E-o]���g��yo.�a.�,=�"���	`3�O��+� �I@�?f�U;U�"�CV|U\�߾h��B�klB�X����FӦ�*�TC�"�FCC�^f��(�Ass+��$87����7����Z }��ţ2:������Ǭ��7�1a��}�����d�����Y[�7�5�H�;nҤ.	$8�1k���G>�~�p�����h���&�[o���r��x�#H�a�S���UH؊�9��� G���(���<t5hX��+���˘4����������w=�p��
�9����q�A{b�/���1-,Z�Ʃ�>�J�d��L� �0 ���gD=͵L�ؤ��f:�MJ.Fq��� �O�G���rA��FƆatt�~H�����#~�k����s2^y�U/p��h�"�Ɠ���d�u¹:Q'�m��Ieh`$���?'�v:V� Ǟ}-rz�uM(�y��."Z���L�g�zn��X;�����'s6��s����ːp�E�`Ū!D����i���J���3�a��v�H2���bB[3TX��מz���D��7�� �|�����mM������<�S6G� ���^W�>5��=)�M*�*\&� ���%L����]��ƪ��[���&�p��Gaz�P��K���������x��r����c	{�^p�KP�n��pl ���a��?YRw?�u�8�5(-�ΛL�Y?���~��ƕw<�o�44���7�&
��[�20��x]`_�����}��u��x��w�Ӽ.\�˽%���}�)���Z8j�-q�a��H������'���G�X;��(���4A�o����̪)	e�%��z����U0�:Ț���߲�EW�;�jޠ�L���;�[�mT�բ��}�{�$��!|��,�z'|�[AOFG�����DzW���ev�c^���4L��IѡW4�9�F�ZWE���kp<�Jb��#�P?"�4���c+��V3��>�`��.������s�c�@}�+4��
��!�]H�}UM�E���I@����R6ᔋ�8[Nz��9��Dv�>��i6�*��68�@,Z��/�LbNɅ�q�shk��<&�U;�f��#�5�r@��:����J��eL�ID0P�a�Ր��Tj#�U���b�ζ�g�����1�\j?DxQ������g�~
�5���n>/�)����9A��;��q�k���& 8vM�@�@Ⱦ_��2;_�b�d�,�J�h\�M���q(�g���T4��ch�_H"a)����tJ2'��9��/G<8:��م�V"�L���E@��w���'^W+`��g���%��E�����s���7	ir��fT�0��}mۑ�#�#���QI*�I���l� �X")��T��ګ1�{*��Sx������_щ�t�Md��j�XF0�Ӈ}�����ڂE!�}���(�ư͎;�S/ğ~�'��qNb��%�^���;֭Fm8�H}���%#8�WOaȮC9���q���kpʔ��<��+X���+B/���#!-�	�1h[ԫ�;hh�Î;m�w�~Uw���at4!�j_#�m�kH�F���X���:%(ٳ��캐ӹ2TcE�6����?{�n0�X]�hL��$�8�4��m�\�c~qbM�x��O��{`d�:<���8��1k�mq׃o`Co
��Eg�����PN���6�a���l����J������ba�E��;4���N,]ׇ#I1g�����'+6��0F.�y�e W���b�¿�
Q�����D���"
�Nɲ���Dj��]��ͪ%��H�4��� ](!!y5Ф��tE�#�/�oX��X>�F�ۛ@�����i��L��z�F%Շ�BKV��ҹ<6��P�55�0Y4U��ɛ(��g�1�Uѐq�P?���|�B�=�pNj� �g�����@F�p��� K5�72����bL��#i�G�(�aGH�V��+��Z�*����޼����٪�.{bVΫ��3� ������5z�r�[6��6<�~�`�B(�Ɣ�Z���Od���"�n���mV9�Z5r^,Ϝ�Y8��i=C�T�΀��j�*
�d���A%:ǅ�b�(�4�0�a��E���v[L��;n���z<��_p�G`��X�3�W�[%�jI_3�!Yѡ��Pe� ��^d]Y~�:Z�ꊨ6*�]g��؊k��c�Ѕ�����_A�I���'p���W��~�V��Z�G�~1_A�Fe��J@�n�jE��UE8B�<9ZI�	a���������L����QG}aK�MGFg8_L@"x�fYT�HƲ,��E�#l�7��Zf�U��+������ܟ�(�:����Q*��%�
�E�:Ĺ�'	Zv�u3{c\.�����Z	pGè������s.��KiU#~&���Rg,Yz�l�,Q6�g����\�xӵ$�M$F��LIQE�"�N�V,��u\(z�U�؛w<�uIq;�'r9���
�N��r%i��K�GR]*�=6��=��3���FG{��a�m��I�_�{��&4ơ)��x��?�'�=��Lq�h���ݥc����b�n@�~�ݥX�̧x�f��E�I��E莍�S���ǌ:c��'@�<�w��9l)�����r-���̤�.|��G�j���{�U^:&J��{n�Λ�}�����͔`�*�'MA��a��`M���Q;X�E0�Y�#�M ��6���D�D����\��ɢ��SԆ*|2n#�9i8�4h:��9q�켵It�c#�6��
��,9r�����
G���A��Rf��5�(;B�".8�"�v	 6-K+�,L��X�ҸN�2UEY���0�"�
�ĨGOl�P
G����v^Z2&bpuj��3�xqP�Y	^\P?
T;����u:""��쳒HY���&��+�s���v�^�[DZ(B�¡���C3�r0u�+��G.�Y~^)�T���w�^^ά�b8#��n-,n�"l)uh��aU��ɱTK��U�Ja��Sm��N���e�{	��$��=�XVHX���ϝ�r�7yF6��m�A0ɨl)�7���[(܇)|KSaV,�jE�%$��KӬIX�b]�������%ne�����*۰��mh�n���@�3�:��x��e&�Θ�[�{!�n������w�~�׸��[Q�ԁ'��7?�1�v��v"g:�|B|cf��ps9(�j|��)A	�P���/E�j"��l1��W�*��\�ע.d�L�^�64	d�:��lZłnSl��]�-�H�=s�`����� Be���d�k"�07^x猽���/������]۲vݲn��7����Qҏ$� ��2��ᨂ�Yƕ�Tc��"��W"�+�+�d
�;�aɲ%�e�]�r�J$ǒ"�@_��R%-�O�!E��X���A��O�{�6�-�iBr�av�@�w@�W�ohC1���T�M{�2��04�P�_�y�\Ti8�Rэ�2�-*����#~_&o"�_P�,���\�N��30����x$�o�H�e�㢮�c##8����?8,�ן.[;Ѐ���/��������X�J�#�i뙸���Q��d_�19�����p���G�@sC\&������8��}ѳ�_���	DCx��~���Ǒ�ۨH�,P�烤��]f���6��m:0,Nv��5x�Ϸ"ѷ��y#�RN�.f(e3'��F�p������|�ESS3^{�51��+U�V�X�B!����(���V���b������\��l���}~rN:�x,�9��5P�c�"ub�i�-Oc�R��w4��m)���\��z��_Ma�����duA.؎��0ܸ��g�U`��� ���&����5=�5�c;�����t�d�I�}'���>8"W�EX��ng�4N֒�����es��_�_Og�[��q�N�UI�b��n:_����T
�o�7��~ųSƈH�"�i\n:[
��D&Q��k��8v�q�q�V��,$.~&�\����,:��n�VU�N��P����A?33h��Yz���f��q*JN@U,�8��Xf��Ҽ��o����{{���E�����������r��yϏ�֥}�c�#.�8�6ّ�L�Ha-:t���Ǡ��բw̖�0�j�����VgE�:����+�g�!OO��TT+PḺ��Y9R�9(V�X/.>� �d�V讅�꼟}�E���ߣ���|;m� �>p/,�%Z���H��[A|�L��w��q͍P�0��H �&t �+��u�0��Qt�@+� _��t�b)��Q�=2�g齢��J���U���?���I	#G�=�.�۴�q�0Z��w��p@�R��Pd�~���/�j%���o�������{����;w�-�f�m�O͓I��dCpea����c�v��]C)��vY.A$s�f�}�b�-�����9O�WP����kU=�y�*�3.��%�,6�te���5?f�����Ds� ���a�L¯:Hm@9�BM4 ��Ac�K�s.�t�+�LJ��C�̘��F'��������6-Y�H��1��w� �&��B�c�IfV%��JU|���:p�x�/O�qBrJ)7��3�C�Qf���Yn?���9����&��]*Uƾ�԰,<c^}s��:Z��{���=����DЯ#���� Aw�y
z�xQ��G"�'1��sd���R�N��K|���F9�w�`��O��Z'2��PX�����mZ�|�t��l��D� �G>�2���D�!j���IL�6� �����n����Ladh���Md�
�P�H+z�iA��ȢdÀ/�Yt��j`���1a!Z��ĳ��ϊ��[�����y����jQ��� Oq����dBʶ������*mbKH4茥 hj���}y�euu���}s�CWw���@3���1�F5Ѩ!Q5&�F��Y�q���������4�<wWu�o�����>�[Mc�?��o-j-V��U��������&#Z2x��0��:�G x����Ql�uL
%���Ҳ��Lo&��uj5�;��0���*~_���ǒ
�7$�Z}�Kq�b�tB�)�*��rr���<��d��td�c�%)�9U��K>ND�=ϟS�JScҴHcAc��$V��4	�H��*�#5�|�܉Gp�9Y�0�%�l�L4 AK'ɖ�E a����g������c������� ��K���涯GF3!�1���/�ū ��.Nxd�F�qn H$z h]F$��qމ�M�fD���F�6�U�G�B,hi�$��d��[������bNuJ}˝/Y��Ǚ�����֯{K�,W���.z;~w���"<���M�!��ض`Z��-$*7���8l��_|�Xy�Ѱ��mS��Bf�`�mX�z�蚍4pዳ\ �HJ�]�q80,��K�d�C��,�Lw+
���D~�4`q�/V0�u0�h�p��$5,Q���o��k�^P��������#�k~�\*�Ƒ��В�QLCS��������b|�D*�.��4I,M<'6~��@75��@8�%�7/�c��T HN@�1��%	C��a���~rÝظk^�,u1y�1;ׄ�� "�v���|Q?�*J6U�@��ٹo{���8aږ!��E#h�f�	�����S�3^Gjf:�0B�M_qC��"��?}��\�f؄k��ٽqwd�p4[��|�%����o~[v�EhT�u("+հs�.��*b�1a�"\Ɲ��H��03[���B�Z�.2�頕�^�Ѣ?{Eǆś��k�7����h�waJ�4�F�����r�cd�t����,��8��d ��1���fn5��~���'m�5�?`wͽ9�G���o�������,��l�(�˒����?5��N}���;�؆��Bq�!h�%���*��KȘ*WR��
M��0֐Yed�����P��j'�0�9�$�(�� ��
��'�̇mӏ��$B��}���aM?�L�sԓ+�F<���	[X��լ�Ҩ2�\� 4m&Tt/�ih��f�8��a��O%u)�5���5���>�qn�����=y�� 䚁�E�9�FCgA�
2HK�������^\l���,�c�	S�Tqb����z��g|�'Tf�v&E�&�Ȇ�5�;����&���b��0GA����<��uXY�XՄ�u'/�*TE��2���Or������7!�!*�<Q�5�̦.��w����U2Zrm@��<��N\⸂��N��L-�a��LO#\�z*eMP�qe3͖��7B�D�!�L�>"��?�<R�M���E���$��{��ۈ��3xũ�q�9��W�\��;�nƆm��k���g�]Y�o	|����32�� �L����;/X��-k��&�<�4���7⦵۱q/z`̈�T�u�����1IL��S!����׭��l�7��z����%�Q�-���t^�ԐuۢC��t˃ϕ������W������ł�_� h>11}e�R:1��N��� �D$E���hzF���{�($��}�խ���i�떩�L�B��"'q�yi�g���tH�v���,B�ꩮ�Z!Jc�4'��qfk0L>�:��=����Ә4x	=I�>�N����:z�)�X:�;m~eGGxhym�aq5_HX��-�7��9316�D��a����D�U�&�!��Z�:�,]�+>�a٧�ڱC<��u�z3s�B�b��(����s��a�	9�p����Emh1Xر{N��(��ʥ)cr�Dw�!	*S���Q�~�[�d#�|xm�J.��fH�DH�$���C������&"?c����$�*�EG��&Z�#����+�����������հr�rLO���]��e!/�}���Ci^�Gf�.F�K�����6��ig�B[*�R��޼o��oq��o����}캾�    IDAT_��k�(b��=k�J�Y���	"6�- �(1��Y/=��Y�tѓ�j�0f�\��K��u�Q�@%@pC�-r#�11�	q�	�PM��I���N�S\�Cچ]4��*8���'i����pG�K��l�l��I^�E�DT,Upl�"wT$yq��-��|>�>�H����38F&p��	����d��]�F�Я3d�T�}�)^,W�u>�D�"'Y���@���@V\;�@*�H#���*��?�P��<��2$�3�+U�
�2ecl�tOKR�\�����4�z65�B���z������@��n��ah�Î���
Ic��g�\��P�5�h6:���G��"���.w�q�!�~�
�f�"9�D�*��??ب*�:N��������Q,�gp��8�����_ބ�zI�a��n�s�Ix��߇������Ǻ	am)Z��pkЌ�8G���񁷬B0�߸��8�ԗb�N�͏��ƽ#�5M������°4�%�=7���>�\�7�����b��_o�ʯ��}�x�˖����+?�9ν�|�y�R<��v�캛���~7
i�o��{t�8g�Z4d��!�fns/�ն��g�|��t<�[8;;�h�!��uY�eFQٶ�
��aYF]׍z��4N#�6C=K�$�
q�٦e9�i�Q:��B3�c�uĉ��,E=M�9 �I5�) �&*�B���L7k1�a�ڳ08İ�%��F{Q����<z�DA�c��$
�?�!���G���W-�K�PH[�X��:Z�i�H�hS{M��RI&�C����������c�cӮYL�3$V�=!ځ�B4x(j���)M�{���p�`;�9֡�@h�yK"I�X��Q)����N��6�RAh���e��t��TC��BH�xb#�[.��� �xк��|_�x�-����BȊ]UL4��P7,SA�~
��'��-f1��� /Xh��N��/zhOl�HO	5[Cw����^��){\�P���L�A ���3'w6S<��=�����S���ݨ�k70�`?D3Z����m�YuI�>��j	Ydt]!��(K�f���a�5�%1�k&]Iڄ);P�fbkL�#Id�"��+�'�YOq5l̎���Ų5ca�-	�`%TT�Ȅ����FI���MR����d�Ȗ��⾚DJ�@)S6�i<"w���UMp��d&�q���*�K�%3�yϿ���焝&��X5�+����W�lM+
߅Pi�ϓ�h���\���j�B#�A^cY��@)��*R<��Ґ�g\�-�ٓ�g��(��~��緜+0��Е�Y������������?������0h��5��)e���$�`��U0����0�Pl�x��˜����Yܱ2b3��k��f��W����@�{C��T��D>6�lB��6|����S�P߿K���ϟ����:,X��W�����/\��P��[f�ן�	���X�{�ԑ����ˎ�񒕃���?���G�|�"q��7=}0�2ںrUag(vk�&�Í� �F�b0���y,.=�R����7���3N?�!�)��;���<�޻[��ް�� @��B<z�8��S��/ޅ{��w�G
�UP�8�(����ɵx�+^=�bA�W`bbbH�j�4�u]�(
˚x���0Ija�����V-�n�)O4f�Ovs?�=�ܜ����뭖f�ͭT��C��/W���|l߾�5��'�/�M��а�m�^������le��@��\-T��̄��Qd�Q}
_x�F�؇Uˆ��٘���l�c*�������#�:vAG��{r���<�~/v���k.;�X:nj�è��b]�*ҀlXS��,�e��c^��8S�������2��z���E���}�x�8Hh�\�FdŽ�e�#�߷"_v���Y���j��;E!,R��L��K�T�8u�Si'Vr5K�庰H�!ɦ�`#j�$�l���]�=�����vZ	ki��o�T)���b�:/훗7v���B���=�4&� �����l]�51��t<Ah�k��\ӻT<�QY�&WZ��݋��.$��څ����-�M+D۰�0F�iK��,w?5�,&b���d��`�5.�aIF���0�O{+��Y��T1'r3qSY�j⥯�����yu9�q�$�= ���g*ŔΝl=�w�,�,RR���@(Kʜ�ſ����|�$�67�����*���@��kdp�!��'?_�؄��0� �s5�,p �r������Z�_ϧp�>���~�HW�9{*��߆.� �k�����'@B�)�M�)IRc8���P��<(���]�"����% _!����1Ix,�*T�l�&�5N�-�	�4}1Ѩt�,)TP�&fA�;g3"�zІk��m��#1Jd�IM!�e�S�h�"P��;.�Y�����4�,�I}��v��߀��48�F�����?����,\8*3��;�E3)`"���6�9���G"�]a��ܪ�:���q�HF�*���8���z/�F[W�"��+�+¦��U�VO��c��v�����
�l�mq)���������O��6�
�����׏��M��_^��܍K��f���/�]� ��+wb�T�N�S�Y2��w�X���=�g/Z���:��<�ח��{xVa�Dc�?}���Z�*0��nق�{�,B�%�Ӣ��8>������Z�[p�a�%�����)���:MNl�L�����P�*ap�"<�~+���.<��n<�q?|��]b\' �=D�nRx�%K���n��Bl���('��4�b2�cK�e$��$�[u��s]�b��8{��03�A�g �ȓ.^�%��4�����p_+�-7���Dx܍���q�A���;a?�@���S�kBxSV�Lf�%��[E	���h�M��f죯faf��^>�3���[`D)*.-#=���v��!U�]��Xȓ}�ex��ڥ/\��cJ�σ8�$�o���2���>7���{p%ڨ�0���{��d�
�0˽�����,�	�n��{�ֻ
�e5	waH6QqNx$nr������U�� e[Q���eE���D�f��T��ߑ*�E�X��8����V��$E�b���-�nA�Q����zNu�5db���@d�D|4S& ��R���Blc�a�|��D�s&� 13�SG�(�9'inZB���di��Q6edb�Ë���RqZ���!���͑�'�<I�R��n���u~7�a���J*c�����I�d���)c���b����[�D-RH5,��y�ZFBԌ��jr���KkE�v����U串6�aX��2K]�} �?CyH�8���3��b�&`K/b��i��ה&�����3H�j����(��N��!����|i�g�����l�v`�&��{�+�&,��L6��])c$!�B<�#�F�1>r٥x�Q����p�wJ���%k���^��(��ލ��^�Q�Q�B�����}�$���=�M�ZC�Q3�ܑ�W��&�C#A@����4EI�U�"�fP�,�z����?>�q>����ߺ�[xd�V|�{�b��U�ߊn��K_�r�u��֏oƻ.%��߷�ŗ�{��(|7CD&/�H�NUDX�y����:��x}�_������}(�75r������_��^�37��O�˚�ә[�[��܇.�1�*���5'c|��ǟz
����{�v�'�`�:ʅ.����L�)�x�E��������������k�B�D3�!���}wdڷ�)\�BEٰh���A�_IRa>���MC�\Fk����!�A���]#:0Q��AHG��o��S@Z4�5;��SU�r�THzd��f#���z))������6�.VF�|:�F�w��*K$!Y[YIj����Ӱ���	x�9�b�����W��?�q������;ox�k�ފ�_�r��ݗ����y�c�������*�/��n\{�-�pϽw�_>�7��/~�'�܆�~����|��{��~w=����Kw��SBDrIi�-�P�Z��h�'��"���D�H9�8ܟG)�6U�Y2N�חύŌ#9'Uh�C�ۥ@�� ��btc��a��F�_�?�Y4+�}�؋��팚|I؄�p�ͦ���
L���"b����c�d�w�*�#f�e=D��3�t��NV4�������Xv�)�<�Sa�0�"WɀǷb.A�.��<��9)ʵP����Y���WE��?DS�A��y&	z����=GG�Wc��وR�G>
]��F��׬T0E�G�`�%"/���8�B%���22�{s�]@XY/�f�!"�?4i~yMSE�S�>E�B��Q5Ll|��5c�\VszXs��}8��,s<���I#��ߊ9���d� !�O
2U�BU�'"e���ˑ y�(T�;���0E�����3�g'�����<�F&����IP 	���tPH���J��!���y��Ex��6w���X�V����C��� �׈C@Fo�x�Y1��$��v8V�B�$v�t-�i�j��ȼ����̗T�r��g|���|�[���; ���o:s	�����op���>�L@�q�z�&-smu}�uwa��A�ia(����鵄�^P/��y9<oz��gNz�~�s�k��9a��25�Q���oC�_������̮�8��S�Z]غw/43��m��D�Иe��ʢ>8�N>�Ttwwab���3����S��ظ�[gf7Ҵ��(I<�u��qJD�d��JNl�r��B��*�D��@�H�LG�Zٳ��j���s4X%��(�<��7;�V0a��r�3ǒ=z��O�[�J�([bA�و"6)�V��<��0�ށ��G������0`k�0��+$*`XB=���)�^�v�㑻ŗ��9���a\|�e8�q��o����!���~�k���W���u^����_� 7�n~t��p�>���,.{���W����_"LZx�ފ�׮Ǉ?u��b8Cˠ�5�>��Q>Q�o̧F����E��>�q��	*&\�!Y�)4�C����t�p��X\����GO���T�ƛX��XŒw34="H]��@!��4D��WG�G3��Zu1�[�Tcۧ�0�.�z�O�0���9�XFC�y�_O2��9At".�.$=�J<���F�'lḩT��g���9y���?{3h2RQ��2���<(�!�q�0�y������:�u1�S�=g��H~�F�)	���]A�C�����b:!��77��\�^�Eڌ�E&J��M�O¦T�n���<�M���Q����g��Kr��@�|M�
�*���#"󁆢4��6@�B!�y�-�Y+���>%��+_�6lI��}�>������� �?�AR�.Zr��<�>o��}�X�a��GJ&G9W�M�X���/�{�R���ВfD�������S*U8媄5���qKS�s0dc����Y�=�T.Q_�[���w��.���Gc��߻�A�C�h�SR䘝^�A0�#W���T�&���o�'�|�!Ʀ�`�X}����?���Ȍ�:�t�v�S�j��`�k�ej��_ >W�=��������w�J�z}�XП���tfF��4s�[���/wj����[5P5h�G������'���s��Ė�ę����L��T'ƓO> ozN���&�]D���.�ꕇ�\+brr���_ⱝ:��AKE�<�NԄ	'r�u����r�0Rq1`P%*�Q���Q�!�9�S�f��2OҼ�P�`���ª�b|��t���v�+��.j�#ԣSM�5V�$(�N_W9�Ri�	[�1�&u1�!	=�)�����7�}:�N��/ݺ=K��ͮp+&V�T�g�VDAAd��;x��;�]���Bl߲�j��v�ݽ��2ݮ{j#F�"S��훰j��暨7���Eb�M�u���>|��B�(�-B0�x`�F�и��%@����HHj�5�$�q��ɩ'4�V�t�YF2�/]Rŧ�{NX�}�)<�uL���o�W|���N؆U��!��ª��b��u8~�q8��c�ο�!_�G6����g�>�-]�u�s�:`�/Aw���0�3�Y�kyC�1�i��ɽ�X�����aIZ�K��[�hs��k�י2�g��g�~��t����q�sڼE�|�Aa&����ݟ[�r~4hX�'�LO)h�XЩK'r�����)�н�[�^Џ����<]o#(� `0�^��ҍ�S&�w|=��(�-��<Ҟ���$�Y�8�8��Q]U����H��_�k9/ӥnޑ�c�Lg��9��}���	�Ӌ�O7ܻq?��]��{Y�AQȑl�؄�T�:""�3��j&�\�����@2�{�Bt�&��c"��i��i0
lX���- yS���	'�I����I�2�6�B�`Aw4���r�č�h蕌��]���N�f4�3�����4t���~��96�7��x���5��q��7�9;-�i�M��%	�"��r��۷��SE��v�܆���ŋ���gX
}��Bt/�o������a���&kʙV���N��'n����__@��}(���;65�y��o��WY��z�fK
zJ�s���~XA��ß��U8��Lozqc�W���	L5�1=���h���4J��Y�B�O�P�����q����w�o���"�����Va��4R�<!J��3[&+�b��i�q"����L1�ی�lHRi��vh��.�!v�ZlBwm%)�d���M�=S�OJz����^ƻnGע��e/%�}�L)��Θ>ќ����jS��*	))�Sa�sĵʄpC���S�e)ؑg�C?�6��2�h�bg떸k��`#�Iƣ+���h�R�maG�ԧ�?;)CC���j�`�k.2�){11"�g5'��Ӂ��m�����5�t�2e('��2�k͐r�2��܅�0Eh]��´-��QA:�����z�)�N�-�ad�r�J��:<q�o������4�#�x�Eo���al|�KG��
��Y��7��W��
O>r?���wqܫ^�5��|d=��!��
��wٱ��E虯3�y
#��W̰j���@Aj⁵[1֢1NI�r�ș����@��\���;�ര�8',����d��".аlϟ%��z@A��F.�~����i��xX�+p� QQ��I�+p	߁itP�ZX�t!�	��ɏq�`��pݺm���G{��Ǧ��
I��HM��&k1sc��U(�Tr���'����_�����W���mqݟƢJ�3�@8�O����%�k��:d�� �(�X~�#��P&S�,}��ș�9�`�>_rm�
L40
P�2�X/�^:��o������|ڴ���ԩ��)2信~��̒�@��l�x!Z�H� r7L�DB5��R�#$���j��Y�B*9 �$���������.�%|���p�i�p�M7����{�k�n4gp4�BI��e��0S�B��`�5�jo�FGa��}8j��b���S�ȒQ\�oqʟ�z�����o�� �V��,N�v\��W��C����{�7�-c���?n�ī.�t���F͢+�'�d�r����9�7�>��/<����uY� ={��B��B�U��S(�Q,v��w-FWAy�O%1����=�MSD�e_A��m"���吤\��5E���eNWL]72,�t�����(31�d.�X�U�B�h{�z��C>��m���ӎ��G�BԙAϒa�ܵ�C� ��J'�>?����)�Q��#>���H�'9.L`G���e�L$�IE���:�2�/�"(��P+�����lcRք�K$щ��+���ȡ����|�e!h�P���x�$j�,VfA�� 1ۈ%҉���((#3"`ʔ*]���M��0���Ot6]DJ��N����P&�ĭ��$>�+p�Y�����24���a��7�{o�P��\��E��է��jm)v��aG�P�����ßŅ/?���;���������ѯ� �n܅�YZ���I�9��E��'    IDAT��}$�J��5��b�3�~�=�z��p6~|��G�L�N���gn�J�xN
�"�<���@����8��--nO�v�y�]���t�T|M�%gw�D̀�U9��8j��b1Bo6�W�K��������8��'waS�@X�!��b�#�8�P�b~� s��:C	Y��W�ă&o1�Q��c�� `�H����+@�ET���.�k��1�>#��1&Z>vR[Y��~^�L��b�ͷ�uA:����� �Y�w9U[b�v.Jg%W'JЗ��3��G��5��4.x�Y�g�l���WP��rސ��Ժ�ly	�aA���I��PRr�Y��<�����t�J*a4WH�i��[(����>�S�W����1�V���~��_?��o�^����n1��`��LPg�l�"�a�g�nÓ(�]A�H�-�*r���zBb>��eسw;�=�8t/A#(b�c�2�
k�<L��E^6�m���]�B�g/B���L�'ܿ��K�~ӫZ�QdA���Fդ�?z��7�ލpbVt�����	��������¡���vbf�7o��P��`�ɧs�U�@���[�7<��]�B�Z�خ��1���d�&B�xAÂ��ND�"�Y�{'��Ă��L��`#C�P��a��X����=�n�a��m�Lm�mZ�R.�9 ���9e^���◷�
�߾��٬��P���̇���,�,�R�#;�L�2�]����CXV"��{g.s��H����]U�D}|v�a��S�טP�TC{S�"x�E:�b��R��NH�o�M_�Rwf�Z�]%�����(U�j�]�|M8
�Nov>v>`�p�G5q"U,��|K�<��%��<��dTa�o����]p8
���uZq��T�w�O���;�x��&��0:���x�j��oߌ��v��֧#|��?��_z�,�g>��8��o�!g��>��w\��;�N���	GG&��-��x���q�w?��n����_}�+�}��'�w1D��l��,��D=��L�s��P�������ʢ6�v��h�wE�(����T>�{Zz;�Y.���[\��hd�+�t�P�i:a!����O�����5�`���_�,�[s<���>3�����Vi�B����S�ݒ�ı��^�2�yS�@�(���������^�������.��������iЁC��fE�Ϛ!.�Fw:��HH[�吣0_Е�<HN&�o�r�@
:���lL��1_3��8����O�����On���e8��cp�ӛ��sFE'6��-�Y�a�j#��0�Y��O��;S��%m�A�X�8Mx�"Rȕa��c_��� ��ݨy{0Z�p�^���N|�K�AowEx$	S��D�$�140�o���7���O:ݽU\tћ1�`H�T�k&�t"t�.��];pܑ�Q�3\q�G��	��i�y���������<���j�MGo��;�<�ł�B��_Ї��0s�_}��SX��0BH�S�@�qߛ"�9Dp�ۊs�[�����Y5���?��?�ꈣ���/� n��0@__�^����\��G7���}��)g3�}�1>��Ie�M,\��,I}"��g����)���9�"�4�)�D�SDg7�^����ecM�*�l�Lu�w�!]0"�|SVƲ1��Z�S�aE���D���0�U�蜎�@}&�M;�[fQ'�Hȍl�Ȣ�SpE����:p
>
ESX��(���3sgs"{J�1M��:�qR���aT��%A�tu��>5';2�B]y[~�d�ќk��G}=aIÑB��<Xa0S�[-�6�E�;�`l1�aT���%lf1T�R5�\�D�����Ò!��-���G�T@���Ԭ3�qno8j�x�`�
���w?�={'q�M�c��z�F`tдB�~֙	���^�����Oފ{�ނ���kX�7������ll"2y����$r��h��d�_D7P.M���������5\|.�����'f��3�P����S)�J?N��p�k��͉��w�*��Z�����H���=,W��.�3��V�,�s>�f�D8N[\n(OzzL]4�]��4ׂG�S�A�u���x���c.���&�I�������ݰ0�s�̉�^�E.�"Iyc���yAČ}��]�H�r��\#��'����$5��|K!��;iK�B�ƌ2�aIze����,��>��� w�~���MSD5��h��p�嬉�OE\���p�I/Ţ�ǝ�m�l��ȀU��ô�J���D��+�Lx�a%�G�6�d�E�47���UP&k��
���k�殻\���G��W�c�\t�;P���y�譢�n*�������F}�V[�7���/�6	k��R�\�]�keLL���FX�`q{?��l�7^�[����Xsƙ�������]h����[n�ǋ_t�����c�5x熱���ێnV#"�m�	;44�wC�$�$G�,+ן��:>����K+ذ�^���`fj�[@�Z�c1�8D�XǞT��̾ �=:�{֏!���E�{���߰c���DEL�f�ͮ���T�N�n�!5�ZV������gTQ��$����p�1'ഷ\��6�a�~�d�ʈE����6v��p Qº�MlO
HͲ]P��� ɍ����͐�&��@����.F�֊��j�.�:�B�,>4:�P
z6;�4P���G����E�AI��S˪gpʖH�0F���U��a2�h@c���%J��MY�0M�P?�F6pkN~�ĥ�݌S��LF��':"����!�T�F��d�kb+�5ga��gA׈a��+^��1;;�{_�={�a��@�IҐ�g�3�:�\v��{�,�Glv��w��3���aO�B��f���F �BR�h�"��H�Ì�E���eX�N;�k�3<�����G�;6!�^(��Y�uf"v� 'F49*��9��7��T���˼��:��>���N؃���p�"-URY�U��J(٣Ď�@5I��l�{�hLa��Ţݘ�g1���%DY	�Q�,���*�J�����="��bb',\�Λְr��a2�SgO0��"����)\BxD����\(	UV؜�iDX����l��ۍ��$t�ŎIej-1��(_�g�J����Y}6�T��3���`l/C!�aY�8|� V�a|b�g:�=���h��H����c�V0�(	-�i:��<�y�^!Y*%��rg�L�@"M�.�!$�M�]��Jc�{��3~:�>i5���?���7]��Z	��X�d�"�/�عs;������W^y%V,]�CV��嗿���&���F�J3�}}�p���`�3�b��-����ƾ]�P�?����L���#�kw�+ q���%]������V�^�ܟ���۟�w�{~pס��b��P�Mxx��P�M�˒������������ܗ�FI���c��ub�Z��i�F,=�+��O���8���.��!�/�	o!g�y�*!_a��8M�L�(O�S�A8��ӄ�3��
zR&sY�`�;p���l��~�*.�E�N\��3xl���<���A��EǟA�R@'�P��}���j�V��F���2D0mS�4�y�Ҷ*�bd�*�D�ãB?r���K�H��ἱJ�h�j��Up� c�
B?��St���xHFh�K�q� �@/j�]Q�ACٱ��=�n�GR#�mDR��Ly\��$�"!�N\9�)�[E����i���G�<y6�9�8�i�aa�$�Bx0�tu��:�n҂?��xŢ�Đ�]G٥������Ϲ�O�L�>�H]j�c1�IO�
Uh�öB�����ntZ-u�y}D2�"I#QaT,��[J�֊�a�f:E��!D>5��R�L�Q��x+�;�*��V��7Y�(���b��}>2����1�s(���9O\�
�d�E3��R�O��hD�Ч�鄁z��ΖȊŦ��1]h�k¢�h��$Ŋ�<�y�kM2��V�q��������̞}w�D�ݲTz)�R�9�3�^�z�FVa��{N"L��Ơ�|�b��j"&�A����T�~��S��yx%����n��Z�G��aq}�"���0��%1t�>��-i���&9$�C�8�k�O�5H�ba��"� C/�4���Hº�8v~��.��\'Cc�c���/ś�=_�ʷ�{�6<�н�٪㨣�B�1���<���]�������Î�!���n�M���� ��^��%ǟ��Z��[F���%ؾs7�9�Lu�j\�����գ��\V
������C�u4��x�:�KnY��ƿ��C�5�$�udJ7ɂ��Dcv�J⃨�t�m����X���w]�:��z]9�D2�Om��M{�m_7<�v5t��~�܇!/��U>�m��Du�t�� ���uT~7��B��Y���+2�j^(��/�pƱ�������s��;g��~[�Jv��Vy��гQb �4䐊��r74ӕ�_pt����d�4�W]$�&\Nt;�(��Q��h�mi6�jQ�l����o4Q-�ʔf�@�q�d�Ҹ����ꐜ�iݓݢ�Гq3�^�FI��1=)�`���\-"�D"c�4�NO~�A�aMH6r`:Eq��Bnɖ��i}r��
���s���J�zW���P?� G�ŗ:K@�\�l-����$6y����.����.��!+��I�B��PC�n�ʠ�rji"��Z6�(���oe0"�Â�S�Ĝk"#N^����� #���j	S�I̴}x\1�ע�>Mr���ؕ�-�z����"y>���:��y^�;i��n��3�s�2b�*9��������?�8YJ�AKYF���mL�#B�ձtؔt�W��a�>�B���q��b��4���[�|� ���&+f8a�0�ΨMI�as����m.��*�bs����Еb�Δy�|!ҋe-�`���'x��y�;��X�8�/Ͽ6���uH%��MYH�cNR�<�	C��JI��.4�$���td�(Y�(ij��L
�q�IMdC���,ʥ�xf�O͢P��n�b�-:��nH0����#7t��u���p����g׊��޻n�!��΃�T�0eq�f�����w����FKv�<[x�x�,���c�G?�����:��نc�?��g08�e�ō7ވ{v�7�KG`������S���G���ً��"����޷���]��!s��;da#J�E��H��}�4�B�S&���3�.G67=�{��ͭ�<v�D�0�
�;:$e����������ʜ;[�-M��-1o��7�W��%�aBXJ
��2�h�H�����G����(���ul[w�"
���:��gˡ�0���W�	���DZ�]l>;	�2o���ٻ��aTG�Eҽu�[��*��P����������Pvk�b�B\�Ov`[1���sphh���,���?*��n�(ת�� �G[-�CwQ�`�Iz��`�R����mWr�}�SMEt��� TP8�R��:�?�v�Bl�Nk%[��S�Վ����`i[��9��OXB�Ua���Q�c8ެؼ�Y(�d��5wo�=	�u	�9���I�kփ=؍�zFb���̮���'�҂C��
�{1"=�O[`2��aƕ��nH��?Woa�`NB0���xl�3б����6��]�,b|���ØF&"ZCOj�u����i{������8��d��������BL�y�ߡ���2.�,��Bœ
��\Y+����FG���� �h�Y]����涋�i�#a�5*K[v۲"�Yy*DN��ʡq�F"WL.�#E�Y�҈P�g���JV�F*|^̅��l�'ձ��a1�wǩU�
��y��� �����dLȣ���ҡF���'F���'Z�J'��|�=@?>?H�\MG!���ً�k��}��┓O�ͷ܀Z��]���,�]�X��t�1��:���$�Q(��!w@E��f����s������o}O?�0�>� �z�^�	��G��?����$�Q�Ro�	f~�@^FW�&S=Co<��C}��a���X����>��җ�W?�&��x�;>��M��:1�sOZ��՗�s���v���Գ����>r��o�p�\ibɔ���uɃ����֥���Lь;�]rd� � ۹�8}�}�F	��(:R"��H*oBG N�k#D'lIA׳����͐�A*d a+\��-�<��$YI|db�	���Po�0�f,��B���ى��bt����W��_�o��!��n���r�A�%�&Q�ZX1څ�ˇQo���,b�x,9m�A̜s!c��C��>��Y F���=%d+�,ž͓�	�V��׀5v��t;D����1�}e˖-�cOmB[�H������T��8��1��&��0Mt-�oX��ST�$����(Wlq�"S�\���D`�2yE�:jG�X��cع�	Tz��*�oS����#��8n��CVU����~��+�\��MI�[�n4���W-�Q�:�Y9����)fg���ج����X���4'q�Bk�_�ѥ�x|���ǮN1m})o���ג�P)v!i���ۉH�0R��3����\�Gn�	ǟ��������aV@��@��p׮1���ݹm(��c=��AF�8��;�|G�\F;WA$	���Anp��</��������ehT��Ih,���w��H�:�|
����C�	�>���|�̍Nc#Lռ���D.Qk񙟐�:?�r�5M���e�{�<��k3�����T"��T�UYQщO=s�ڼN=c�Ɗg^ԅ���w�n&�?��z@'/���l�t�O��2��y�ς�8DؐΣ��U*	� ����d�����Ed�@ܞ�Y�;ƚ�C�J�듨��G��h3IQ���݅fǇU��3�16�tC�.D�t�厮��֙��V61��!|����M�|)���Cgn<r/L��r7�Ƣ�i6��K'ǩP*�C��4.&��2Z�&�P��I�!��,F�Ȫ�CT�(cff+FG�Rv����%�ثc6ʰ�'y�z��/�r���G
���z����n�!����2-̗I����/ �4��}R��$-;� �c��Em$$��E�w"G0�byI�.rB�< =�.��=�d��$��%j)Bf�u�ӟ/�*��d2q����@4�q��J�d@�e�	}}��	���p�E'bדw`��}^� .�;nG��eO�jg8��עg`��?��[�ށA<�~�����\�ahW@+�D.�4��G��k��w_�c�9
���f|몟��!�J5,;�H<��n��
��ǰ|���%*(�,�_�4'�d7�^s8.��]������^��a���x�1�/�N��迻	��J�l%0G0�g�����X���X�p	J�E\��7��P��թ#K�,�g��ވ�n~������j���Z^���|M|��&���b`E%�+�]�]�ݍuݍW�{�^^;�'?�aր����s�nԺ����b�Ƨ�]�097�2����<�������(�J	?��|���\�ِ{_��B�2*��,��t���vaim��{
v��n���_��5kp�ٯ���܅��<0�vAv23��+�N�F���ǲ֐�lY�r�<�&:�  ��K�r��o�}����hAg�0ϖW�#�ݵ��w��Tx��
�<:+���rx35,
�NZ�O��!1�l ��	gF�i���f�М�Ũ�\;OM��[�'b�L�("S�<Q�:y�IV��Y�"�S����d-���#JB��(��	`;�Hj���ʫ����ԕ�j���#�S�,��CL���DQ�T�'|�i���g�6��X��b�$��f�B!�څ�p��(u��鉇159����_�����=wѵqΫ��˖�緭�?~��F72�h$��xL�2�e�cf��Mx�����W����Q�Tq�m�	ϣ�Z�I>�Bġ�a��[k6�\�A(��Z�"��yGB�\��%k%B���6�N���@    IDATQil^^����)�]�'�U��?�5�z����~���Ю��</�������ȵk���d\r�l��fC�\8�+�Q�V]��kp�O�MD/v[�<�ͤ|ɁU�!��^�Z �hfb"��V�B���M��0��L���mDr�3�K�9A�NS
���Ȯ��R�`+�l"ؖk��4�
�:�G��f|ﳗィ��c��E�P��޽�ɏ���.��F�o^r�[f�:�h�&&���kW�7[�4�j��P�ڂ��)�ͩ��ы_��o�	�>�0�KPEZ��}m�Ӄ�ob�����UĒE+�]������{
+���_�w��Ocbl����[�íw>����J?&&vbd��O_q9��{��{`�����vz	�V����;P	�p�-��U�<]�Ep�>i�X�B2s�G��9�-O<��N={��o��v/
#� hh�t5!�[�fJ(G��p̈�;��!�>�^�ַ��w���⒋^-���V�X)��7^�=O?�7���;�O�pՉ�����L�%˗K-��g����}��È�
ܨ){���0ݑ�t�{����W9�a$�旾�s.|������qԵ*�� 27!Xr7ʐ��w#���[���v˲��VT���9Ԯ>�c�VI���)M~ol{p���<������8���FQ5�t�mG����iE��>�V?�� �k!���F�f�EO�����+�~�:f'lQ+�Ȃ�N�jY�`�S�S�QJJ�l>��w��!�^#~�~Ue�}�_�ا<O|`rɜ����=[П5�Q�u^�&/���z�]9�K�Jg>2�>JN�'�#�E!������<c��"�"��o�ۇ� @:���	|�#�ūNZ�ݛ��\-��]�[-W�������U�M���>�5I9�3s-&?ꈼl�V�F��Mx�YG�3�p9.~��tH�P�����՞k��ʍ�4�"H�R;�Y�7<0���x�e� �Z��"l(܂�����{�[��Ɔ�2���i�������p����8�?�+��{h��m��93g�L��sso
�@���A)RA�"��E���)��J�H�%��z{�~�9���gn���~��.����%�ܹ��o���t}���|���>�N��MW#No&'���t(�
��@��m���Pu��&�C�tv�iJ�cJ��M�1Ti�@��:"�@!c��Q:����7�D�mj*��ٽ����8:]�h�(�Mz�T�!#$M��Wj@L��H@/�3#P�a(����o��ѷr1�2H$U���=p'��*J�2�Mq�Y�A�R���A4��E����a��_�/�xnv?���U�����o����'�{
[m3�[Lm��Z�kbvL�r4-����?�7���
�u�y���q���0�f1֬\�>=����w��}"rMx��'�d�|��̋��ii������[��>�뎸���@5M|��l��6�o�¬�b T����ڈ��AL�����H��Ճ8��Ai�Z ]���P���$�pj4JB��c��m�;nŻ���9\�B����L�)��zb���S7e������2��
"�! @Έf;���Q�b��nL�4	v$���2���U"�P�.vC�(M<�l��eU�*��^B�V��<��<*z}n˺J����EI��<!J9ͺu�ѳ�Y�r;�EBB���G�s��
���� w)F"o�������2/��[  t�ٙ���������#�Ȣ�l��f3B�Y�H�mY�(�8<���y���J6�ld���iz��=2�xV��D�A�.a\[�T}C���(0B�.P���x��!6a}?���Z���ތ"�Q�$A��)��G���xl����5����O���+��FPA�<e�T�Ђ�k���a�?*kF���#=B���\�S�K��#nW�7b�f�w�^��Ǣ�o�k�U����D<�B� r�F{����p�K�`�ZP)[�Y��èT�r�ё�(m+#b��߉+.���<�x̟�&~0�n@c�[$"�=����r2����e�E#(�J�܋H���.��j������6�\�3��q���/ ޺z7v�s�K��ة����W�S�`����;+g~���'G	���?d�������%	�8,R�~�V2F�����ҝ����Q�R�-��QM�$�nś���1�E؉,t-	'�0�~Ǆ���kS~#Rt�]���Z�;7��ى�WWבo�r��,p���!��F&����7]s�&������&��{%�~�y��0G����d6��>L��%���l 8�G7`���E���"
�X��.�*N��ECX�r��vh�4*���ђ��,��on%,�|�t.��&c}��nG���~��8��mP���u˱��b�̷��Ï�ؓ��]�?؍��㚫~���aD,نx��{�}\vݝ�ͯ����)нaR� ;^���H�(�3~,����T3º��)�R8��{PK��fͷCB���U�R�U=���cJ����)ýX�z�<�0���L�k��WWmq`��w�O�3�X<�eT�z��܆�kW#�ڈ�w�&�B��]��
ғ��o	~���O��vl�Z��w�R�;�\�����<8~�Z�j?�J���H(!�B�)wp�l)p�LF�o!D�MKȤ&�,��b�"��.�G$��;�Q�ư�.&��.`Bܤ<K�o���[�����}�ב�s`��θ�3���B���]!GrG.��o�������׎�t�+FM��I�>!��{�QA�q:Ǒc��r ��C��0}\F�Cx��70u��0P����B9���U����ڰ�'��bzB�d�����;% 1�$�)g�tN��e�XA�UAF ����q��HA���̓�D�rM1��	�ҾjP��L@fT�Nr��IAt<!!R�f@�+H�U�K�ع-��r�~�y,|�M�R1��b�XA:��3)�҉[`ֲ.��p�p�t#�:�E��ttQ�T̲D�zf��&�������W���}{6�]����8�A6bo�@Kj���(�6M����H�6�>ұ<\���&Z���/��#�Yׇ���0�4Z���oZ��?|�����g���#%�oz�����-���
�����ʤ������a�.�U�YeRQH�:cG�hV����Y�W�55��P�LZ)��zQ�C_�E�ΟG_8��z~2+�g�H�2.��i�M���v����O��;xڕ�<�CK֜�� N�jZ&�XC�Fg��ԃ��_;eޛ����N��傰As��n�l�XL:�m�����z*R�0n�6�{�58���2��A�����N��=~
⎁�@?�锐��504,�"E��>R��T��,@8Ǆ�[a}���>�_=ٷ��n,[�>��mG�?{.n��fl�����3�����@���]����!A��U�q�o◷?�s�q�9n�6ԳZ4��\����O�������d"�j���4�Fx�����vl�YV�V�
�D�����T�r��)�6)P�0Vv�chhH����{fL�b������ա2�]�뎻B����ܷ���v�h�cʴ��v�4l��θ��3���uH�|��{=��k��ր��=�c�������9�8����8���-1�~T�g��c#��DP%�(0���A�%�ZA\�����#0��$g"�=�
�� ���+f���S���M������+�z�������-�c�<7�U��l:~�����d��׸F9�>/\��VѢ�
�	��A�A��
��q�&i.<N�잉@p�,�ڛR���탸Rz*�0:��v�����|3;
��u^^ч�P�P�iF��A�z�I��$�E�a�3��'w�N��T�{U�U�A���'�O0��8I1h�G��u��E������B���,1��|�P<	��u������wMD<j��Dm �����a�o@upL��t:�P$!�w$B*Gg>�T�;�bX�Ǔ�)�H��È���������R0��1!��#��=�(n��:|n��100���|��;hn��(�9L���[[[�qlذA<	\ז��Ϸ�g�x]����c�m��o-�ٗ��t3�&m��/C�.c"+��)�����:�O{<e�oy�E�.n���D�\���e�BH��^��hSV�7��ah�L4%��u��0~�$<��s8�أQ6*�,�kC��������?��ﾍ��o��5�PƴI�1w�Ft��`n��%��E���>��M
b������P��dX�O�gq)�����$�n�"�9NUC v�VM�W���E��k�F	�X�Df����F�cT�a3^d�|	��xX��!L2\6�r����4��G�W�=�:[��!s�~c��qQSr&�f����`i�K�ki���툻�}�>4{�;�~��T�1o��a�V�0{�l��1�e�5�!ߊ)�:Q+��ctc&L����k��K�#��➛�GC��=���\FZM!�e���)��U@դ�{�p�M�
Ӷ���0.��	�y�*h�[�`SU�1H:�� 2�uw���$��"Ԙ��U��jF�(��!��ߏQm�`�L(�$4�Uc��ZBCs�*SE�� ��P�Z��0
*��}���s�&��s0a���3��~�]1�P��2��1����{��-?I"��@�A���-k��\���a$�H�D�&�*!3��u��D>�#��d��]d�8M!��0X*���c���|�1MݠFO�sG�jԧ�^�f,Az�r"�]v1sa<qDo|�|�R�Y��aD� �b �3~'w%��D����bϠn���?8)��<w"^���Ǖ�~���r�|�1�}���������	炂NԛS��8���M����L`F,]7?�Fv��L�4��ͿgS\m}7�ɝ��U
�)���Q�/�Ӳί�]� JE���ѮTq��/��Y��[g�$�s2��T��'K���ފ��tzt.�
��� J��IC�ќ*S���x�����E8���q�=�����{��/�����b\g��Oz��D"!��������}|�ZD$E*ـ�pE$M��#O8[��}�=�. �H�|;�p!��-����>�����}6��;R���?���<;�@��� ݶ,�#]�
�*� ��q��u��~[��0~�x���X�d1v��nX�ۋ�k6��q�M���U�Y��ʕ�P,Ր�6bݪ.tm��X��{ћn��L�o��Q&Y1�"�4�|���[���D
ah��c��Ν������0!2��Z*�v`W|I?C�EJ��g&6!x%�Z-75�\!�����!8�1:�>�΁��E(و��v�E,��g��2�=w��q��U��SO����&,��ʐ�-�5J�&�B�c;a�q���D�f9<�N�cTk\�Y�{z`jH$�P�O`�h�Q�v�Ԫ}�57c�N�w�Ï4�4<�ݶiG6�b]�jtuu�ԯ�-[PRT�d3T�����D��T%��BOϜ�ps��(�x@�!�-C��p�gA�w	3P� �\-B�&�>L����RL"aE�W	�P�2%"nw!��tZCE����pሆx�	C�׵ul5.�&Ǳd�kyh-������7��Z�y̹g�k�LX�fFl�G"L9�G�%�+bA��v��"��(U$Z�g5ӫ�u<a~s�w�K�&�-�DX�y�Y$��1N8�����_��7R�=qq�naz@��$�p��)>��>����X��E9~��˶�֝I��i^K#=x�<D�2J��B}����b�=�A5������LƜ��k��2.���o*�;���
qa��+���4cCN��N6�e]�Y�-o2b�[��`���҃��%h œ�u����/��G�=��8����K����b����%P�FR�4`���luJ�^"	qD���q���b(�ВM �����v�/�=wߌ�֋?��� zz�1fL�pUʥ��<J�i>��Bgg'�z�������ȑwA�aT6�r�W	cC�0��[`�=F��@)� #>
�Y��+�|�Q�M��mͧ=����}s���<����T<+�f DM�mI^�J#���{%�q�n������G�W�csG>��(�.,]�7g����q���t8���^��ٜ8/�]ۋd�	�P'�u֗\}��X��@���B���%���ƣ��E���o^�%�,f���i�]M&��R�,[�ݡ�,ɐg*:��	AdB85"�)V����)Ӳ�JJ�˰��r�NHR��*�B5ѡ���HB$_�W=	´fY<������S#b�E�j:�A��!�*k��F&��*��d�l"�ێ	D���۱R��3�b�0b��l\+�D(N�W��2�FEI��-kFl��M�k���L�V1%U-D� �p8!�ȋ����$G���Dw[��aǐ��#��
#Z����5��Y�s_�dV���
ٵ1
!pK��Wc�0�Ѯ4)�$��
]��8W"$��#\���ؾ�E[6�����RH�y$ՌX$
�bQv�t�����d�tW�z���:�.�ҵ��Jȗ�&�k�1=�]U��*BQ��S n	v�U�Y��AN+�T0a{Eę�gnhA�	�o4�u��\����#,��sGI�RB�d�N�,@t��VG�V	��%d�2w��6�P�4Bb,�+��G�x�zl�j����gٳ+��t4jaLni�Wӡ�X���!U%7D�tZs�OYk� |����ߜ�?rF�ÿ^Љ.���F���)��z�22�o^�eż��C�� 4F�id�OOJ���U(�~h���['�]�@�w9���bm�d�L���ර��-@,�&kD_ՠ�x�h�}U&�p�G4l"60�j�:�X�w�)8�+�a�g}�C�z>I�^`"à���f����^{���_��:�\!��r~1ю��Y5��|�z�hh�@��qX�;#��s;�4���[�?~�	�����?u����zD�%?����}�W�;��9[�;ACr9"�{��ב��x��S%\~��h�V!b�f�,Z�ېj��|Ū���<N>�@m�����b��r����6f�~��8�����`���Q�հ�Nl��-W_5ތ�/�1f���O��áըK�)aU��3˚� ۛ%�3��������G�0	U�M�q-&��c�%DlZc�ivh&�r0xFg⚪��Q-�ڏiQ(a]�N7�G���M$8y�*����XЍ���!Ӑ�;�XET�D4���TU���e�4d3Y�}Qb�$趎M_*3��#��jQ&B�4l��,I!��3
|N億`x�*"iʗW?�db̨N���A�V51������Ԩ�Ё��PF�_s��%�XY
���Pl n�p����=����#E�m�5�d�tSZ&�ZE�g3�:!�fT2�H�`���:95��kɄ5��͸P���JCHƣ0,F�F-p,H~r�f�����!"#>߼-e�tŋЌ�	d9�#�iK�J��~Nm5���`ژ�8�wc��a���a"F}(��gA��A��W��:��Xw�Y�Q1��ú�b�v$s�D�.ll�"lB���xԢ��cP|!�96�M���4�D]DTW���]�z���G�p_(k�{1�qsi����(j��sV��!(�a�[�A��?��9�>�PKq����t��>@F~���&`�;Po���2���B��QD��;����C�
�bQxM���)�p|$2�8���q�C�CI4!�j���ĵ0�%a�caD,�
��z�s�ux�������гv���P2!��4���	��"���,�=��\��>>���T*�7'Z&	��ڛ�X�|!R*p�Ϯ�Q����/w#�w�՘�`#Z���&�L�2Y��ⵧw����?���Oy�}���?g���<4{R1�)�`��    IDATnzG�*|�*�T�ǚ�Xy-f4Up�%����
b� �G��=C:'l�w�/Ûo��~{��-qo����q(a[tLFY��`��_�@w/N��gxc �y
�%��eWo�u#�������z,H�J"H�2�i���ҢE��Lg� 4"��җۃOJ�L�����u��qd2TuS��e�M�=�����XP�q�	�	��D���|�h��Fq-�Ѕ*ez�ם�<S�J\er�%2@N,�H��b�8RY�S����\�hjjBih��ut;�q�*ð*�F�"I��qDyػ�@��
%�n�P�1}Eē�M3pKQ$�<͂�9��%*
ؼ�/b#�Yq�c-�,����M6m2�h�,�bQ-��+�f�Y$�eK���0��	Z�9���d0&�qR�P�)�+5dY(3���&��r`�-̜?�K�)2}��Q*����_o�� -lA7ʰc	,&����@�82��#}QM��|C��gAg`���JX3ȣb��Uth�0�vX��6mx��g�d�<{�X> ��@�nr��N�^+�J�v���	ĮM��ǃ[���8Édo�P B��e�&.��Jowz���P����H��u�-�@�|���{|�1�E����?mQ�-s��03Q�q���H�x]��S�,6>#�.�WM���0�O�����D_��A�ya��I������P�75Ҵ�u�u�}��\
�#�|Jdɵ	�0[3�Y8]Kq�������D3f�èY�1�ץQ��x���u1x�9�2��-P���$t��F$�Fc&���e8��p�e���+.Ae�]+W¬֤�+���ׄMg�Zŋ/>��^z	�\�|>�v�����.�7m�ƅ�)��1�AP��O=�wN<�<�����w�������]���Q��bF�=�������?�y��G�����������^1����N��'cY7�j�[,��!^Z���M\��}����; Pu6߂��*��5���@6��ba�.pz��6���GOw�
v����8�;?��V8��`�20�W�H�	�Q�B�8>�p���Mw�a:̅�(�gJpTH��p{K�ALK!�J�V��Ɲ,��iR�.7��TH��&��nI�-��k�S�}�I�U�g���C��rj��4߈�����4q�;cJk��G��%�+�|�T�������N���Y
r���C|U�0�iaOA�V��m;m��2Z\�+���&�JM��J?�b�yeX�E�G(�=�m��y�Z%B��&2&�с&p3�J�H���
*�����$��#V��{O�e�����n�5	c��P%��h*�a*�ҀɇN�~��@�b ����\v�sx��w��SN@s2�{��Bj#�H�9��W���G�@���<���ZD�M�E�Hi��\
z��%����^�R2��ƆF�I��YB�~�B��c����4�+�����g��ةx�=}dTI��ա%����6���3G�&#���&H
����JK��;�
Dlۇ�=��"��2$�Q�V��	DBR������<V*�|��bJ蜙	,�A1�k���B��LM)_}*����g�tp�O+Пv���9R�7Mun@@�2�y;A$6���W
:e�\�P����Y�۷g�/N��nX���՘�Q��g(�H�4�"�Es��mw�7��OC"݄x.���	;�A"Ո"X���y|�����n@�4��'�8�8���.�s2�9�_w�ux衇��:��Cq�׾.$9^k����^Akc��Fl�;�L��f�y�������?µ?�'_��q;�b}?�]��_��Ͽs��[~V�?�u����So.�y��l3���e���P	�;:�Z!Nf�+}�NW}� ��yP�n��*;T5G�ZF�4ČE�G���x(�&J�����^J�T����5��ο�K�(&� �oC�M�OǨ`b
;&���@�]���T�gU���
,z�e��`�;�è=���C���r!8�I.�9��E�C�s���R�S�DF���XV*2��<M*x�s�rz�������\�a'��o�e�QC�h*2)�:���rf;?��j�D5m�
�ݾ�,za�!h��]Ln�|B�X��:��2Q��Tj���nH���O��ӣP��Q6�u��`�$�*�	M�l�0q��1g�r�_׋pC�X~<'Z���j0��ޤb긼L�kW�5졒l�ѐ�j����g�<(��眇�� F��0E���{c������`����ݳM)�^ׄ;�����H���vx��N<�q*���=Q҃~�� |�_b�	I�{�	��Յ_x��+�m�����fF�� ��%S+ Hm*�!)�,P��،guh�6�Ԟ���V��~�Ս=�:8v����K~����+��Z�	�,���Y�cpH��oZ��������:tv$�I���RD��㎟P~]jG�(WY�~��h�E/x��3Lc�6�S��:���b�$��� {�؉p�&��k�P�?f�-�7'yVz�䳋��zA�!MP0����c�Ȗ���T�G��X�W�&�r@�����!/���?��eA�8�]=��	?�-(����U�̅�N>��W^p��d
kG�	F#� ��z(��	��_�aH9A��"q8jB��,�nC�/����^sҩf���/�z_��н�Kr�-^ �>sZ���DCC.^"�_��)�UK=��&L��m���R�ᘨZ����y��g��z�q��E��,��^��'}V��3}�������뭥o]��{;��`�kbn�m�5�I�:����1\�����3�rјi����H!��D�F�)���QМ���n�	cg`��������z	���b}-%�Cʹeb�KW���[�C&e[s|׀e���r�,�&�0`,H�X�Q'Q�7BgҔ0ҙ��I���Fb"a����[	���dd���i�O�0$�.��"�H ���aT�EGFA�<�ￍI�hm�bɒE��b�sʔ�����J���è ���~L�Rrq�rM�0���^��2eE�L�B��+O��`X�9GP3�3i�j!�˴Pu�� N �F>�B�(!ݐ�<D����T|/��EdQK�����g��>��6
ǡ�j�e��+^_�KY8��G�����gc��W�燞����mТ�	�Ȟv��p�/��Y�ӹ���Ƃ��"�2:�R_7&O�N�	�p4�'�ÑG��\�m�wL�m�=�h,���l3�W_���ϯ�q���<��B��jJ�Y
�ŝ8�c@a��aDؔ�B���K)�Ù9NS"��!·�b�%Lj���Z���e����β,�K������ȁI��H�s�GoV�C��-S-�Ԍ3e��#��qS�('�D�\����@'�03�k(�*E�p���tƶF&u�-U��%��>�;lw8��Ę2>ק���J������@!�״�k3��,��n���~�-��/�g���n�ȶ��n��`1�B=b��1o|EV�����^&�:	V�ff�#BE �Д��$5� l��0-���<�H���֩;�f��x<[�� ��]$�н�cnsP�B�(l�P�\x4�Y�_��:�����G��^�d(�+�J��)S���y�����Ż����gr������Y<��b�
,Z4_����L#��`V�]�]v��~"�Yha��౹���	[��+���{�lB�����}���̼��E;&GI��W��zM
zX�%���^�]�8��£7�"��*W�O���.l��%��r͕�FLXf�g��{bG�`����/���+8�;�`��Bz̖�,AQ�Lxυu��Ch�v�<$bI�<�Ѯ%��N<Q$Y�P<����Oㄯ~���UĚ��c4�	��N�$(��<2�oR�xa���HRbI��A�iV��KA�=�zZ�.��І5�������~�xD]]�WI�8�-z����+���H[������u!�:IL
��8��
"�$��_r����<�L*װSbB�*Wq+3�r�9A�Q_.袙V�)�\9��Z���1�h2*iP�'L��5}X0%�M�G}�L���9X4����� ��c�I5�=e4����ذ|<�`�'�?�هPn,���Һ�x�������+s�\���k��K�E<BGG;~r�u��'��G␃��W\�m,]��Jc��񷷣�1o�0��8��q��G �����~m=yT{;Mi������1}7���9X=����E�;~�Q�Ӛ��ٙ�n����%�I-*g;wל\i�)��{���VL��l4��X7PĆe/�P���ָ�4P�����fDU/~#Eed��W�RhD�ɴ2v�4m�O�R���½c�L�D�a�\wE$���%s}}�E`9J�4G������ȐL��g��E�^X�������Gx~���F=���e�`��qv�@Ἇ��O��7�6��%�˵�EC]�V�7�b[/�\g�@ OLx�q����	�/@Z��O;I�W^x&F�j�c�\\�����C#�։�B��Ɋ����A��2�ǙNW��񟟎��>���[�����̷a�ݘ�6e�d)�|����koo���X�)���ј�&z�L�W����GU��T�:�m؀BiX.�|�4�0��J`Fcd�SW�����m?��7N跿����?�����AA�U���k��k:���xu �|����|�.��i@!����4t�M�a{6lwH��¾*:^�2�H
�[ḳ.�����£'�K�1<T���J\�B�����z+6,�'���ڮ%�>���䖎c=c'LF	Q�{��xi����q!��Ra٢-�q(Ѱ|�z�i�"S��x��2�Iw\(l@>�5���߀�H���w���݁�&����N��wf���_vU��*�Q�A�g��i�[�RR���Z`V=4�PՇ��Z-�hjj B&�%���r SJ-��H-�����u���a��ֳ�Jh��K�<�T.�'�:������Z��h.VK(5d�-�j�鈅c���`�Z�u+�|b^�߇PbB�2v�����G�(>��C�r���l1�IK�<Zŵ�`�_���w��λ��Ϳ�9:���Ͼ��t�rꗱ�>���܀�*3f�?s_�7,�_�z{�'��e��x��Yh�=r��8�qե�A_��y��x���p�a��<<�����߾@&�G��5~��y���o@55��/?�t.#�LFxL^πu���i��Q&�
e��hť@P���t��Mh�J����4q�$Afb���X�ǹ�	�O���Vv�#7+*�T�Y�=N�#9��uF�Ԧ:#]BT�Q�,��i���p��|~��|8uS�,~I?d���(p��3Hd� "z~^�������t��h3$^;��}�I�4��~�Ԩ��|�|j�?�_�@���Vo�����ػ��(>6�?�n84�?�?wϔ���fP�Q���b����¥g{h~~��h�g���#�%�B˵Ʉ�lM<EC<ـPT��8`/�ѐʹ@���[� g��������(}��e�QN\���D�F�m;(�4S(�"T��T��q]�q-)�6cF����mb������70}�)�X�n�~'��׆��=l��W���S&��*пvϟM�>�Gn{}ɜ<���é��Lj�kPC��SG�4�u��Wb��Y��D��
���fa!���G&/IH�x�M/xƥ��*�
�SI$8�ě��+����&(�`�q�Z��qh�Al��q���Y:��s���Q5���������A���)|�p�|�z���G�y�}C�$2Bl�2��"Sa��HS�:xBm���f�3���.!�f_/��&q�>����wa��p�7��}��Ͽ�,��Ы�V'ԧ�r�QR��UD#�0R};.�Jĕ��;[��h�g�2�4|��f-�	R�|��aq kln�QP��� ��6�FCS�@p�DT��M_,��ˎ�{[{JzC�*�vv��K.C�\��/�6j.ι��������÷1������?�J�e���}�����Vz0�$2��k>���>��Z���z+n�ͯ1�=��x��٘���hՌ�|
�=1�'N�g�-;r(Z2��ko����o�~G��\c'�t>�w�1���c��p�Bt��5k�aT�k��;�}�0��6O�|Ȍҟ�Y�
�L�\w�n�D0V� j�E�=�Y�wK+��4��c;�h���	�?�K �#�n�a���ؤJA@�K�@���������_�#?�Dx�#V����w��ɇ�|�F}�2��'��1��Y�-@e�J [��H�_'����>����Z$J�D�q0ɛ�Fp�P�Ai��y|�!'���\���ҵ�cj��?�o2�٬A���~G��w�Z���$�xŏX�'t�QB=�hf��Ÿ����W�����[�4j�LO��ʥ!D�8tOE��%37BS�<�e����O��T2��Ԉ��F����W��˾u��,Y�Th75�̻�T9#��p*Y���1|'@x�'/�*r.!e������B稉��Qq\���(%�af�
7��֍��W�>a������볂��=v��̺���rBg�h�"ӹ�P�m lU�KP���s{ۏ� B:��a$�,�U�)�BŚ��e��{���i�T�ea�';&�և�G��S-���Q�}�~(���:�r�H�j�l��ٿ
���Ӷ@�� ��v�_��v���0���-���I�܀W�Z�ED����0/؆gؒ�N�B�D���Ç_ؑ����� f���� �b��)��D,{�q�8�g�|����x��g��%J��pX<�%�RI��I��4
�Aѵǔ,����6Ӆt#�M���ЅbM,T3�8��"�ƶ�V��9����E�C���(:X�������I�k���r�7t	˾eT������!L�0���*�;\��2��Q���z��v��bVtt4�:�e�lm�����4��K0���l�<�w�}���k1�-�u�6�80��1��ؔ�kK�������G�K�)���I�t4�M�q�3�m����Q8��0c��p��64-�b��(`���E$A�-F�z���7�5h�gu��a�.<I��l�
O
:�d!�G��
,?eϽ��X���B-����	�P�ɓ�T�A'�6-gI��9��V��g�n1v�e���&8ݞ�v�������B�*��x>ɧ�����!�M&�G��M��%�:��z���x�,���0��Q6��u�8й�=�ʥh�#M#�N$O��!q�>�SAh���Q<�X|����7ۡs}"�x���R��	��@B72��Q<>a+@���"yA��x�5nX��,����ݳ�A��W�<�7琈�ᇢ0�� ���NX��
g�_�D��pB�1�n��6�*�0�!��$�u�%����a���݅��Va�ر"���&��
%��LV�w�'����l�Ԩprt�F�!/S:ɾ!��jE"���Րn����v���g��k��H�-<��ūN���+���=V��NA�����^��锭y<�*U(���g���eP$Zw��m��.c��_9�1,r��9�%�jU&��de7I��hd�r����;%)R*�������
+҈H<%�'T{��J/���#7q��f�_<��#�H�u����� -�A]E�!����yg��<	����P"�HQ�8G9����;EL٘�V�5ա�@��I8��]�
�s��J�q���]�v�ډӎ?sߚ�~y��VY`Ǔ�GBe��)MV�� ��2��Fl1n����5�X��1��M,S�����^�b��J{Ѹ
װrj��J2\Z_vݼ���$�dR��suʂ]�f�xH4���y�����H��@8�C��s����kpB��    IDATƩg��.��5
{g)�tF&����i�O�Z�r��CS58}+1���|ֻx�w�˿�-���`_7�����Ϸ��ϯ�Ņ�?�c�:�=bg�K����G>7�����pōwa��BGg�r深͌=�jX�x�{��X�b%n���[�Q�Bb���&x�����K��GR��#���,NG ُ�FW5��	2��g+����Y�L�hGh�C(�%Ǚ�>w�A����қ�z��KY6y,�aʳ3���HW�#�E��0���0�K<������|�]�i��A�Sf^����$�Q��3����#�z�_���RF2i]�/~��"GI#��A3�ʧ����������k3��~�����͏4�Ws�Tg�o��M��5�f*��o�|w>B��ϐ�f"'���s�m����^�ӽ��T6��;n��8	�Q1�!�5�O�������d��Ga�P�,�d���(B�,�7X�>\x��8n�]��+/��u˱߾�cŲ�(��v�jĩ8p�ݾ�W%y�׎�`�R�ӱ�N�	ӐU�OIbby���
��1X.�s�����x����W�2mO���8>1���N����w}V�?����?���?}k�,�.��e(ܡ;&<J�lS
�Z����rئ�G�Z@5$��/[�DRC��i�0
�*�4�$m���nc<\�t#�D~}�+Psca:a466���]���j��2,-���wV-� >�0�A��u֐j�D~�t<��ҹV�+�z��[k)(i.S��dX�-2�n�z�a�;����'��]C���}aW�[+�����틨��s��Y*��e��(��Zoml@O�:��,B"����0t�����B�4�|5�6��
���bY�P��
�>��%�C*�F��E�\���H��2a��a7�l6�tkV�]�TBE"�Ak�X�a�ٸ}���kp,�
S�h(C:��UW]�1����m�cμ�8���q�7����V�G�H'���M14H�P����0��K�r�,<�����?AC6�j�=�V!�bⶻ��+~�V�0��ם}0���184 ��X������c��҉c�?^v�@��'t��LL�ֈo}�^��Z��6C��W�Fi�Q�������uu�^9Q2U�)�$�@����oO�z�.�J �u��DX�"���P���(~�(Mq6cC�ϖ�ͧ���ǿ�9]}�ɢ4P^Hq�E�D\w��.�iN�����u�L���.��8Ǒ�J�aa)��
D�B�C/(�����P����(�ؼK��'?b���fc�p�t>B@4�|"��*���$�X\�#^�uo��#쓦����a��L��3yY�_WAd��#�K֮���U�d��i�dZ	"a��޵�zV��ӿ�&u�]u1Z3��46�b���5�M!��5��
|�H4�M��k)��2P�M�ܷ9�p�Ix:�>����0�'��3�I&`ٲ%M�5$b�L���^777�<�)kD�H�e�dsNC�\FTkD:�,ּkׯ��-۱�����>����n4�����(�cj���c?<y�_i�������)�[��'�x|�����=�y蔿��
��(c��*| =@¿�B�r�U{�m^Ǟ8焽��s�b��_><�wޛ�>v�k�{�̙5?�ޕ��ʫx��'�����\k3y�I�[��p�/��m�����JK.u�w �l݁}'���E1�@�!���	K�����K���5�!5zk��a'ݍ �L���
W�����C�E�zUyH2�D����wsE�k=���q̭ ���¯���یϣm���ʫ��ڟ�2u��4	l�)�g`G�%�3�G��'���p�ᇣ���{����8���g�G2���3��[o�UW�/����\%,�o�}�{�9�X��\���v��p�����o�g��{�����_x/?�N>�+?m
���}X�zN<���	�\���yYo:����$I{PP	۲:9��/㤣����ո����s�_�=hG5� �xY��Q1����)���x����ﶻq��7"����c�����i���/��
v�ak��콐���pE�J��x}�*ء4�fw�7��SN��g�p�?���~�?c�z�p+�0Ӿ��г߃��O�5X��<	�#<ڤzP�F�s
Ua�T(����M Y��o>�/)�Ѱئ�a�i�)ς]��� P̼w]�	Y�@�/��QѤ�U��S�����.�A7������o�Η�-4t�B�{���L�aq�yf��0���F�:��}8����k��"�b���,'�^�P@!����
˺��9LdFnk���!iN�����D6O��A F���7�N��l�.�>Qþ��������'M}'�^ж�a5���9�'H1�
~�x��)!��k8�6�N��Bh���>n����h�o݇?�S|���
hniCo���Z+�mw=�[�~^�J.�D����i��S���P�u�$�V���ਃv�%������Q������,�:��t���ZZZdo�&����QW�?���cP�I,]����e�����g��G��/ׄѓ��@مU-�ǽ~߅G������w}V�?嵥��OΝ����%F���b��@��e"�Xp)�2<DJ�[���:����ᵧĪ�KEw��s��-�܂/�zV�ވ���	|��?D��.�r�M8��c�kjƣ��L�T�F���)�Qg�ʧ4/_���<��^~�I!ڸ~
�]X�t)��7N�b*����ۦ�e5Y)��S�G���'a�p+&��@�ją������~�v�&�I�탋�S�V��NmI\��г���=%����܊'��0h�e$�!�k����K���n�r��|:���&���v���O�ŋcҤ�x���q��g�駟���_��n�	˖.Ǿ����N���?`�I08�/��G�(��ҫ�k�1��8���Ï��������{�'�zGq^y�E����_E��){A�畊䚚0P����=��yW|�K�����87��y��څ�h�K�Q��pcR��[v$c=��V���~�澅��{���
�0{�I�i/+��<��|w?:�?�@\z�t<��K�.`�ϰ����H�I4�EsS'�r	�G�Ɓ����aŚU8�KG��{BU�Om�u��=��0��?�B,�@�0<$�4�$�9�Ͱ�HfT G󶊃x,(>&C�D��|(R��e��٤8�8�Px��xOV!���o|͹k��t���mH&���%{��0E�ʇ�'N�ax��0��]����{��U��⟵�j�N��$3i����IW���  E,G��G9EEУ��*� E	��@h!��:��m�����ϻ�@�w���=������I&�����}���)��cdi�tB�>?/N��O�n@���L��(^ӵx$���O$�������Y�j�ؕ
�TF
���]O"p=ˆI�|�M�$�D�<L!�`�W9��"�:M\�����L���}H$#>NN�Ώ;���Os�q�{��Do��8q��Kc@�E�j����_�ӂ@P���uIX�u]�	o������$�|#%X�6�}��W�^�'�x�3�	--!7LE.m��|u������|	�	�e�x�,\��� ��
C%ͨ�f��}�
~��յ���[�%9W�^��	m­��RW��*N�--�"G�� J� .*����&M�A���"6�[P2�P��ȹ
-��G�pJ�����c��J���w�����獲���\��֥;f�%څ0C�jh%BU�����ԇC�Ʊp���pJ��{���8�����_ށK.�,6lى;�?��mذv�O8��Q�Ј��2�3��6�>���V�g'��@F�����}�0�,�Y�)���m���`f[�H�\B"�D_����{��-U��uTc&��C�J���ÃD��"%Kp��mI���#�v(]S�:jD&].�[d�`zp�!3pҁ���Q�,��k��]�v���a����q�m�~�|���b��ob��'�t:::�[����Z:m���R�;w.n��6y�.��tww㥗^����BWW��ڢĥ0��_�'�x�v��+�}�ٸ�{ĉ��������ù�+�s���ݕ�=��%��n�g�Z����X�`���'�=w݋�iӱ���-�V�.���╡�R�O��VB��,�������B������7�#��5;�H�j&�$��m(Z1t�ŐJ'��d6��Б�f`
ȚI�z�W�2����:|��Ϡ�{&M����}g^p6~�����Bh��E�X�r���\��4�L(�D�3����]���z�hL#a��7�5�FQ����L��QW���}��ː��`��*��h�][��d7>��E��H���&v�QHHT�"W:=�_C`�)F�PSYi,<��D� � yͅn����s�0����	^��S�
@�)��Ƕ����E�G*S'!w1�wP��N�.�;���0��e����Y��.!0t^t�u��a�5�ruhFE��Ѓc3��;d���b��/�`����ՈOd��F���� X�߯���@�]
(���<���K�������k�>���)��1",�B0���=���s������<|���HP_[��X4;1���s�=�:e>���6�2���^����i�4CBo���yF=v�_�3N>��nF~`-�}�e�������CH�S����9��$�	1��P�td(Et��6&����dFG��G&ی)S�a٫/¨k��0s���I�Le�X%9w���_}�G������W}X��~A�����?|i��w�.�܋R�]�tZ����q�t&0%�`b0ϩX��q�ǎ������܋���s��+��έ����O�S?���ז�Ŏ�*J�V<��jl+��[�&�"��}|銳�O��P_ʣ��v���^��o	�44�4����A��~b"��ba�N��H46���Hd�a)�(��6b�Xž�G���˳8�C����ը��7��́��K*�V#�pŉ�0�-��	|���a�����ĺ���1���$�@'A�A\d��o���kv�K�,�W��<�����q�wTƉ����wߕ�{�9���n�"F�~=�".��2<��#8��c��3���/��%�'�h���e˖a��b[W7���/?����V�%q��C&�>&�'�)r��׾{�7|�<���`��C#�p��P��c�RE�LM�"S)5�Y)z�����E�%g/��5�pi��Ç�7%^Z�]��2��S����.4O�"Tu���N�`8�S��AM�ҝ˱�'��\���â�������ԋ�E������'�$i�u��4�i!Maj�k�mAU�0���(b�l|�=�>�u�؞Ú]�S-�1@s�6j�8L��C �	Ӳ�ۭ�sn�}���||��i��9���9���Z�_�	�bI	��=�x0uV�(�)���v6���T� Gt�4���W#GDzz�9�%������5�F�c��.���h:o[���
	u	��0b���Kb@ef�`;�誫L2��Tk�WBi�uz(���r%H��*,�����#kܸJɫ"�z��΋	#/2����v��y���	q@�5/~�ض��d�^�أݻ��n���"�	�� ���&��	��uo���*���P����
�ʶm[P�-������{b�}��ek�[��bX�>/NS_��l`��Ů �P1�ۇ�Y�����x���G���O�kh�%�JUVt,��̘>o����۱�~�ᵥ��yc3���L&#�W����p��L���9S0\(�e�ȶ����7a�£�nԒ��ܖ��K�q���7����a�?zz՚�_�2���
:'t	"��R��t�Q�1�GN�b߉:2�
����PFC}�l=�re�(!n$d�4�G����E�����㰍v<��J�,��5t�Qu�zn����&�!ُ���bʕ���_�U+^�l���E�+��k5��Is�l� �Jq1p�b*|�D�����jBU	_:!F���[�J"���}��t�w�U�PWL�H	���ہ����3�9�G~�@�F����}o����&�C�ErU�zP}][qݵ_º�6��G��3O_�#�9Z�����ᡇ�	����_�3f�bUq����ɧ�]��n�:6m؈|���<�g!��3_|�x��%8꘣��K/����Ý���v�I'bú��<u
�{�Y���aptL
g��M���O������阦�X�%խ!��n�^sq����矓b$hƿ��
b�{#�8�3R�	�:2i�F�ju���8ᘃpЂ9�m�n�$�~�-~2U˫FpB��P��u/&���f�U���,��EKC�;�`\t�L�D >w���Έǘ ���.��N�pƝ���ԯ��؅!t���_��dR�K�bgY���p�&ĳ�ٲ�����x\��P����]�|"�z�G�+��)y$\#b1e�K
	c~aD��*N~A�5t�1cp*Eq6,W��,T:��eĹ7�sȍbz��QS�ʨ�Z�z��&8:}��6��e&?W��d�=^���$/Ԡ�q�SW�)Xy��a�J��Z'�_�?ހ������ ����Ǥ�p����1l�1��ר��o��eDS���	�w�s��H���8���v'ȍ�������3i�j�j���&r��CO���_�jH]"��bA��E(8H������[��3���DC}�v�himB%_��9{"�B|�g��_��~:|SE��B`U�dŴ'�U��4>~�����K��{����[��(��#��!Y�4��Ze,m���G1aB+����w|/���h�8�rA~?:E���PT��'q����ދ�N9�w���~�S.�[�C䷇�j~�O_>���ު�_�nN��xB_�×���g&I&u��W@h�j݂[�#�����
=0�"\��l*)u���.�d�$֯�{l߅�'�˗�����hjï~�v~�]v�bHC�Qyqg�=��	'ކ�m+08@�4`��I��7��:Ͽ�z���2C�*�'�B5ю��V(t�b�3eZ�鶐�+(�1�] *�˩��L�G+��T�:�Ѓ=s>f5:�g�$�`�6�|�&���e��� &v�⻢ٵF��ކK.�ߺ�۲�&��_�9N�MMM2��'�����Ǻ��q�z����q���U�\���^ê�k�T߀O9/��4��c����ȣX�plۼs��ųO=-���]=���������\��k��ݵ+�>eJdY��PM��d��	'~����Ǟx��`G���ۈ�9	Z}ML�.b�~H0t6��40cr��b�;:Hb�	%ԐΒ�U��e[�t!�!7�TZG�M�S5��:�r��P�Y��&U�ō��!{�>����_BǜExm� rz,��f���=�)�"�N�v\�M����2�������+u��ϝ��EϽc�6D��Z � M_X�N3���Ǥ�sj�A��J&P�6T��Y����ː��h�y�0(�h��*����+X�փH)̝1U�C�D9ȏڿ��.�u�ذm�b�Mx���	PϚ�Z��o8 c~0U�ZC�B%�~���P:���6��=.�!����Г�+��#��q͆ӿu�&�:,Y�c"�DJ^Au�&8hV־�$�oZ���b��ҵET��)@F�L骫H<-�|�M렦�Ľ��nJ���+m�����#O��k�5/���k�Ώ˜�WB���j��b,�3Q��3d!S�arЇϝ~ �ob֤&,��0lݶϿ�4�3)��b,}�ml+��ݝ�XV��wB�uŝ���9PU�S���يs?�?n��+p�U����>tm�(23��)M㚎�3/rj^}�ox###�_~�g0u�t��r����hl�G]�3��    IDAT:�P�mq�on�| ,��}�8����fNC�vpДĻ�}����K��w�������~��kn]�s:5�L�
�"�*�x����s��8x��ESꐮ@s�/�B?�Q���d�h�¢��:��̲�K�4*�\MdO5���?��lA>�"�j��sgYBX-� s44�,>���yV��,�c��(�m�6��a���u8a��P[��D��4�E>L�`r%j	Dr�t5���Iw�11caAg��� ��p��R	2�+���v\|�"���p_(�$�>�~��o���c�(�Ւ!�$�έ����:�z�)����p�a8����#M�=�݋�3g�裏ƫ��*g��׾�5�؇����o
$}�g�/���%2���O��w�-_��iLo��;�#���%���/���/�k6���k�H'�ͦ��{����t���?��ښQ����SO�c�^���w�Ȋ��NxZ&��ŉCg.{"�j���!QG�" ԧ��<IZ#[��!�`0Jv,�����
PS��%1�.���K�Ill'.9q:N:rOX�(�ϙ�{��w��ET�)pb�(���Xv}�"-ܩk0k�B	�1��Ʊ���'��o�G,�V�؅��T��D�$E�iE��T�t��Y�%�2�B�&�h�΂�	O&��!w�{22yGn�
z��u�8�۷�+`������S�Ō�S�ھ/μ�Y�h��x��qǽ��_=�g_܄����������;�܄3/���k�G�a�e>%|M�l8Bq(�zABف��Xˍ�y�k��P�B���~�����o_E]s'>{�w�iD�˛�	SP��f�������7݈��M8��#0y�!X��0��,��,���nXsL��ЪD��?�����#(�+���m�����_k�IjcP���G���g��	�w5����_��*��K+���bHV�ؿM������/C�+�� �u�}�a�?m&V�_�|R���*}~ #VZʄ�T{bn�p�����:\|�~���Sq���b�Mع�=���r�<K_}===hkk�%�\$�ӦM��M����Jz"�6v-��i+͕W�oS'O��Y��V��O]�	9�����8p�XQm@%���I�[��'������w��������'�Y��e�s#�ZT�Cfw�eh�T�PN�&�0�]
�߷	�S�B8����0Q�i]�#O�n��ߵ$W�+Բk#�4	jr"^{g3
���| +�	Oo@��Ṡ�a��H'�Ѭ�8naV<�l}��G�լ!������G���BY�P��~[�Xz�X���DN�1K�SUc><g��r�<��F64�ST��������Y&~}�������c��Jndw�vF)Q��#���$���8�����o~'��qt�x�w�1oڸQ�_LN���;!�{�WX���8+V��n��SN�7��|�_Ď;d�ɯ%���<w����w�)��m۶I�j�*�=wz�n�^{�;�\x�%ز}V�y�]D}]ZYAHc�,>�<\����֊7���p���`����7ލͥ&���P�dB��q?�������>3F���TI���͘�\���,b��6p~�j������e��vBc��*�T��T1����s0c��>r�1��Ǐ�5cȅm�I��p�p�Z� ���]�jJ�bw��F1cr���*屩{�1�>���̬*�֨�P�KG22�9���b���Ly؛F�v1< �ڥ�/CMd*���&��ԇCfNľ�)L�8X4;���v���e��j ����ҏ�[V�˯Ċw�cݺa44�`ۦ�1�-��?�F���
��K��w�&�_��Eq�R�kIm�*�q$�q�'�=Y��"�e|�Y�oZ�_}��hmi�G�8��D<�v@1EkDPô�������/��[�^�i�\�d�,,ym]en�N�h�*�z��/'�@s�(�Γ�O	���׷h���8�����>>ы���6���ވ����������4"HN�_���Ƥ���-���z��8�P!]g��K��:�D�bc�E�o+6����)mT+�B�(
^J�dkx�<u!>w���-�adp�_~ٔ�3�8���'�<�B� Β<"�����KO��XVdyL^W�m[�H�pKTM���6`��)������^��}�����t#���}�ם���_�A��|�0��=�b�mKw�ɂN!�S��΂�@+��Gqp{OM�����E:A�IWd�E'�{ل�y5߅F����*
�6�3bS� ~��r���(�2�1/<?E���su�%C||A��V�EKR����V�$����\s-R,��a���!�г��pj
~R�<3nHV��p��Bc��JIPA��x5�K}����=�Q����6c~s��n�2��f\qѹh�H��^}|	~w�](���4i�����A\��ϋ�kC]=V��R4�$��_��ktN^��~�0�Ix�$�-��/O,��?,Ŝ_���g?���կ⮻������%�~�m\p��?>^|�E������g>#F�����k����X�a3<� ��{����hiL	��f8a\�����k�Cw�쟉i<��-���Í�xNf&�x:-�^��F�R�(Kz|�3fZ�U؅f4`~G.?������~�;�NU��b��}���9f��O]�-���`����2��(�l�yGL����U�3�=��Gw<��"�fj@�!D'�����C��YMcd���0�Y�:��t�#�o��b�0�@I�R&*���d���!����(@-̧�Rv$�mM��>cz<{�j	�w�t��	�CC��ܑ���5��ه����:����c�o�d�&`���.vu��)Ì��;g?hz3֬^��C7s�������q�����N�"����nr|�Y�I��<u柳���0}�8��n ���܍��o��S���/~Q���%��f;V���m�Y���S�q����c�U��Ϟ�1l��-T�f��4�SS�%��̀;t"����LE��� �i�M�Oh�V���OG7��?��^@�<��\��\����yQU
���%���_�"y�-X�P����FD9Q)��NG,��>����(��&T-ˏa��$�eP�UB��[�D��]�d��:\v�޸�'�_�
}��г}+���yi�'�����G����8�ӄDKw7�Aq�'�P(əB5K���Ҭ�1�m2h K���kŽ2�܎YG���V+
���.Y������'�0���������Y��=P�m®۠P*CKKJ���Hz>���8��f|��Ð���/쒽/�{��s_�ΠX(G�f���T]#r��Z7Z�e���O� E8�s_�]��l�MH�/�VE�)��}���g�ҘA�\,A7R��)dZ;�hl��ШX����,��'���_�q6l��M��$k��#�^���]E�,@G�
`��F]a��������Ơ�u��;��x�^\p�E��EKk'~s���a���:��e�o���5���a�	y�
��4&<�	�����Lvµ��B���>�z���r9�P����n��;�֭[�g̙3G��͛�"��`ڔ����c���86"���l�ϛ�s.��l��-�q�������eK{t<����E�D�r	VeH�+k�W�����x��W
(�ť�,©G����[�wႋ>-?7�1:<�3�8�|�j$R�Xۋ��|k�|d�g��a�	�CY{q��S�G<� R�Ky 4a�-P\B������Ӯ���f����e�p�T'ܸϯ��y�Q
����1���u]��Q��֩�P<I����pqSsp�Yɾ�/07Q\x�yQh�J^�[�ջ',�����t�.x�����ȴ6!�؄��(�X 5f#�0����(p�HsM����.�G1k���Oŧ�����c�\ɒQ�bHIʞD���'�E���.01�wꌐU�6T=w��X0s�T�2zs6�V1Z�-��9T7@CRŤ6�MIt���P��Q7�$ӝ5�YL㊋s9ms�����h�-M�j�@��E~�b��(
������q	Z��G���q�_��5."��ǹV�l�q��,��E�<tG���1�M�t�"��N��kh��JC��wA���6�B�S��^F ����2�O��n�cӐۆ����+/<?��O12:��/���l�RA^�L������yAeK]c��ㆇF� �^R;�1<�/gDn`�l3&L����7aB#e��68�B�0���~�ޓ����>d�����o?��-ϭ�p�����OA6݀��n ���9��sP+���8u��[�;��CK�4,Ǔ�eѮ���S%W@��#!aJ�#E��cvnvq������8����Fn}')� �#������NGп����*d�;hi���E�3�k��l:)E,�iF<ۂ���E�%�8U�CX��ȶTGӛ}��Lb��$oxޢ#������ o)hK'��؅E������U_����Z44���Ǟ�U�R�`��X���=�ooF�\B��`$����Ɇ�%��f��M���/�8�hp���ܨ��i����P5�	Snd~�NQ|�)AcN:�B�$�n�JF2�Jl��(2	�����A��tCŔ=�c���x�ȕ�8��O��e~u�=��v ny;v�$R���H73�b�K`ҵ�d�w㾎�nJ��X�w ����'����Dy����Xe��A�����^����5Tl?���z�SHw�F9n"4����t.l��5��m�t�����(�í`Z���i�[�܏��xǞz>&.<�.ۂ!�F�DX�1����P�8\�Dh�@7�.P�<���Ř��Ý�<*�$��mwz4�K2KD�c!�l��"Id�é��ނ�����yi�ң��?G��#c�Еu	�2�
q86!Ts����sga��0tUθ�r�(�s7ގe]@��}���:+	��!��[A�+��i�̍T,��Q�.i^v	�PA�Q�u��ц:-��2q.�@c��cD��1K!�bQ=b f*���:W#4�^�$��񉂑�&��<���w؋Bv�Ip�x0�������j��nֻ�{������㱶5` ��}Ĩv���,0_
��/��bR��wıGK]�6����U���:��%Z|ާ��èTE�hi8v���&oyG �/\|2~���c,7�o��ĉѽsZ[��W)��gSii<(#j�LDѩ$ݲ������^o7���FT>/�`,W@�u�<�t���ՐGu��<���O�[���?��	��O���O�\�×wLϥ'"ef����S�FMv���i��p��$n��h(#��PFx���h���t媋�HF<���)Il�
#���Đi���m]|)V�݅O\�#tŦ�o����õm�AL�cK-	���CP|m�� }�*��:1T�~˃�(ϖ&�qB�U?�ą!��'�R�љ�+�p҂�oZ�eO�	�����뱽�`�n�Az^������kn��"�?9��:�����9>n���9}��O�=�'|硑���gC�3��r/B|��H��.�'	I,�,�
�:�ȓ9� �H���nt�iDŁ�
�ɦ���lF
>�rX�͕�b�C�+s�i^��R��ylZ�Z�{����w!��qxl�R�O�O���vQI�B#i��H���Ô3��u%��h���Ѝzl�2 �_'�*0��8��o
�?h��|�߯E�2����m[?�8�t�����Z�^���,y�&#�3?����yj�${���Z��](�����A�HTKػ>�W�X�G��^zg=�z4�|��t-
��A%�-+6�.�����ѐ�TE~(����eA�]�4I��ZA�O�4E,e�`E���;�_�h`צȨ�)��)A�q�t��~�[U���r����ϚBD��� ~���-�ެ�S��ܙhhj��`k�]���|�������s������1�i�<uDqx���Ej�ߝ�h"iSa�4������w�B�0i�>�, %n�$�;J�2��� h	xݰPq��ȬI&�0�(?"�RYݠ�D���|������qX����}��\����u�u�=�o����"�G�eN�]�s�DBA�]}h��M�� Ǣ쭄���Su��%��%/�����^?K^[�R�^<?�DN�n(�s�S��B��Y�n]��O]�k/_��.=G"����x-���<ad�1iB��h	��	��
E9?����jKl�M��,��2�#dRi}$L	��ü��D�҈��$�K��o����t����g��<��0L����u�.�5u�l6q%7���]B��#�2ۂ6���R������F�w�`!�gP�cP�&�6���* �!��Ò�`�H�:06���ş��O����t7F���N�[-B�$�U�H�-�C4U�B%DHY�xo�Bb�}�5r�2��%���G��Ŋr�X��m�E�N^ܭ)UĵP��,��!�p�������/���0k\s㷱n���7[p��+U��،�\	���>�w}�*���~�������ؾ�ý��+cBPi�0*�������`l6$"�g��&$(�rYn�� 	���T\U�R���������m��ˣ��At�,�bC}�eK�''�B��D]�r��1q�r��%1�7���>Ă2R:0}�D,:�p��2����a��~��^/�I�$c>���t�9b���<�;V��疼�C�8�>v��̧:2>S�z0��u�u��@��l�lc#�G*�����G�Ö�~L�{��<�Ʋ(1�+�@,���;Q*�,�4�HʜtA�$��:I��wW�r �z������������cϿ�����%�'	[�֥�ѫ��;e80���a��[d���aAX|�?PY��� F�cnD��N��+ô�P�v�C��˗�yӚ0�u#~��{�n�Hc�A�f9�A�n@U�
�T�2���7� DK�$w�YX�k_��ϰ�[�9iJ$x���TI\�8��E��+Gֲ��
Q��L��W�4#��x;.��i�į�Ά�dU�CB����e�d�G}��χ��X]�r��IL�x��r;��	�gN�����z��g���^��B���R�F�Ժ��q���.�E+�ȭ��r�[�Iv���U��W�أQ�i;����F�g��t|d_�y�
���-/�F4D�(��p�wh;��04��"�`f��G�������Ƅ��عs',����.$��.�2)��xN(<�H���s���1R쨊$��ߺj �ϡ�`\A�/�����aǞ��;�|�lC+,���	j��7�;韭�}8������ӫ6��jW':�1�UA̷�%�^��R
yh����q�p����
��Z1p��U��NƊ��x�������ٍ�_����b��7Џ)��b�{U��J���j|��?Aj:��)rǝ"���ݳ��	�ʣ����@���L\PG:]��m��*��3ʵ\�N�c"�&?D\1�sJf3`���6ǅR�!Z�l�5����+�&��� ,]��A
�u�l����HXy�Uz�����ئ7��C����V4��q�{U�u�>ba"���5�U��k�!�"�0M�g̉�25ˈەB򠆊m�����B�ɜ7\kS��֭rE
����:rB�,���V=K&F�����
EI �i�_�ѻ7�GҌ�ŧ��*���s�ʺ!��	P2i��┣E���Ê�)�5��V��G���9s���x��7���G*SkۻhW�8��ðGG#�����Kd$MnB�T̞�7�R�o��[Ħ	�y&Jf6'��+��@�a\�g(5�!��9@��0$7�W���YLj�¶�03M��U@WO��"v�Z�D!1��I4(/N\����� 6�n:K1ߎȕ��d��Gq�2I
�>�S�%�RR���n���Gau����-��>{
�}�)<��C��LZ=�    IDAT�c����:r�¼�t�����T
$V6b$7��B^Tǝv:�:_��v������?���,�HS�XY�;Ej��r6n�� )T<�#/t�֓�XP�1�͡ˬE�e���Y�Y��v��?Bxc�!�:�tȋ��ꄪ���BZS�ܨsUNO~J�jIh�g��,��oB[�m���
$%Fe�!z��9'� 5���<XiRx�k�$����$���=U�B�BLL�8z^�V-�[�����z"�i���+b�L�^���������`[�襨Z��2j{x�ۊ?��z<��#X��
lxoI�b�U���9���GǄ[CB�e���]z�>���A[[���Ջ�n"d�k�pQό�}��}�G������������{v�#S3�g�y^��������O���'�z:G�YDsh�P�t^�A���T�^؁s����:1��!m�Z�߄�[KX�|'�{F��޳���E9��%�;汱�j#V�5�����X��F|��?�;y_�ciБib
����%a����w�������'�p����x<��g����s�d/E�3'F�Z4�3"_e0��V���r�@�t���l�A�ˣ#��~�o���J�@%�3R�]*u�r�����Nԕv☽��3�<�u�.�!�Q�a�H	'ub�:�v���S��W���,�'!3�ˣT(��CR��b�nB�#�-*К�|���t���NB,P�����E�J�&�ʊ��::�"��b��i�ub'�TF����v�T;�DVޔ����4�y��+�hM���S����?}&�ێ�V�7Նўn�ߑ�ه-�U���m=��+W��#?����F#����������x˻+��fĸ�-&rG;j2�c$�8��w3��.PTz�.�$�JdM4%�w00L�ڨV���I��I\�A)/�'cr�Y6't~��4r�$2h�} ���MV� ��*������#Nv7WQ�(f4űwg߽����q�����!+��r��ΎirRߜ��Ǔt�22ȏ��\�Xe%/���m��sp�Mwc��Q�u��4\��j �k�P��o=���=s45K3Br ����2��d�+5E����s�)5�A�H�עk��/z<x�OY�k�6b�lh	Z �o����g#@Z\��"��*0�0Z|����%���n���G�~������@-"��}���߸� I�k�zq(a6���#�n˵GH�TL�}��MmE�Z��L��v�-��/��O�u͘�(9O�A�2�X�lyq����&,>f��u����	?���hl�@���[��/��cWH��z��N轾�.r��-A��sR�	��!�g�)�|�߾����o��[<��*d;�DŨ��ؿE-?}�����z�pB�;/Go&���o{���5��֘�:�~�9��Qڹ
�9�1?��ehI�:���>v�)8�ȣ���7Q�XH�28d�"�^���0��"fv�Ւ���d�s��g��u?���i����p⢽P���{�~d��p�g���;-��dQ:S�Rw�ݸ˸��  �٧��0��:��B��^���B��}�y�g$�X�ʈ�*��:���(�J�d�1�`��
L�UT��G��-1��k�{0�>�� ,@ӿt�CLseB&�HSU�]��WJea�W�Q7͢K�v�WKZ�ELc��d�B�I<S_'b��zsC#JՊvN��{&���[�L�_{��"������9��1���ց
Vn/`�M �2�4a(�G���^��8Q:���`Tǁ�0��FgK!Y�^yv�c,_�5֋O�t .:�045��p�_p&��	-m�������[7~���y?x�U<����������0�k�kte�5��}(M 	�y�qc�`d� ڢs6��Z�t�c�C�|�����>�\\N�qh)aGH�,�P�V+����..d|nj�~DŒt0>\�L^cf�)�}.u�,�����K�9o=��� f������݂�3f��o�#U���"�"����I��֏��QL�܁IulھZK���Ơ?�{�uT�8��SQ%PLY�B�DNl䞱��?"i,�ZsI$HX��pF�
E`��	�PӰ�*0�Ia�S�{Q��Y$��<�j̅'�NF�f9��'���)���w=�bvEe��E�.ֳ�*��e�{�Jm���Ul�A��%lD\�t��9�	]�H�|<�g�{��#"�4A�cn��@���ܜd���*�2��h`��Y2��)�B�0ɞA˒�]�	�J	��	�0�n3���,\u�"<t�_p�Y'cxp CC��0hS�F��|	��!���!
������i�y�Ud3���y�hj��+|���ζ^��#$�H",�a��}�'G�?�ۇ��_<������XHw�!�*d�
�;T��h^�C�p�G���]�E4'M�+>v��y3��/�r�m5L$�c�{f��� �DJ�2{�w�w6��/����X�m:<3��e�й{ �ۅ�n�	�L��W}��QJ��.�S���G��$���&�������!dHe��$�k*b!�.a`@�D�pqQ�	�{'��$�I�A��l,�Uj�]h�
�R�Đ��g�jmF�54�%�wQ-�d�f>�fFŹR*ɡ΂n�	�>f��IF�0�(�7�CO�j2�y��#NI�)�\>��ىU��g������WK�x%��Ld>��#�Ks3�m�2Ǫ6��3�Ci�� �WK�bK�BR�+���`�)�܋����_E�+��9WuQ��pm�o\�M��h�T1�tp���h6|�ZS�M��Ukq����K��w K����am<��Z['\f>;�8��6^Q�'E��p��s��:��*L#-�H�k4���y�'����O���Qȥ<��81dWȞ�O,����'$Z��š&H��T^���6�v�p�,���uE�aX7u�nCx�+���1�Qʏ�*ԠձQ�9����O�z����aG������g_�1������W��Gw�~���7���♗�đ'��o�^|�j�L��KeUES%��G�J��ڵ�5w��$+�(\��p%LKhHs�c"��f�{�3�xW�p�hM�̆��7^�,�!��[Z��L�ӅC�)�;�
c��={\��Z!�O��ؠ�"P#��ؼ�[��Vc4�
�F�߭��?�t� �Z��Qq���<R<Z`���׀Ǭ���Wd�N�D%W�J���*gO��&�C��p���a4�1T�ȖU3i���!���0hn4�!V��3��sF+fϞ-͒��%�:�&�V���YV���X.�ȴ���6�PVzt�L�Zd�!U�W^Ǧ�
Ԧv�R�(�4aR�V����*˿v꟨�G�?��gy<�C���7޽�О7�$���7�䆢�3!lU	��n�u��z���N��h���T)"�٘3w6��g�m�9� 8~ ǫ �q��CG[vm߅��"6l���]y$���c+�à���LK^tK6���u���2,�1j��l/"�L$I�Y��b���yo@.�E���k�됽+�M�A�qBg��qh�'$��t�4-I2jv��<x+��)�S�'!tޤ�4�Eĝ2T��<;�.S�jI��эE��*ֵ4�����?�D!�����/���$�Y��FԖ�y�A��y���H���K#f������Ȣ��FLC2F�A���DV���O 4�(��(^S��H�s ͑��\��������������P|�A��8[�um�����SRhj��-�fܿ��;�ڝ�XЄ�a2��L�>�����E�T08lak�_o���N�c(d�c0�;l2�1$L����לGB�@QI~#��2���ZBIŠ&�v��ŔiG���Y�"����fa��RZ���L����u��;E���G�h�4!pUtoْ�P��_s
�*�wa��8N��';;`Go	aB���P��7���[tٮ'���yM�亀����$� I&�9#H�"�r��+6��HFf�݇6%�ܝW����n���j><7"z��I��I&m�+�
t�n��J�1�T�p��,�a�n��;_,�Q���+��4��e�4� yp	6��d��U�
��R��h���@>�*���G�R-"�1�.ڲ#y't׮"a2W����0���ol~t��߶���L$�.�)B���ad�_�")/$��{,��W�'�Uz15��:E�[��F-?3�:���@��<�1n��(X�4�1դg�8Wҙ����P�`i���X&�Lc3B�c**�~��d`afK6��[g5��ԫ���aA�;�H.nzp��{���ml�U��".R��������c�Iu�{o�O�(�_��P�GEW<2�G��#�� ֙�M�U�FBK"?f#�� ш7��`��H��kDA��&�� zh���3���*d-ŋ�J�}[M���d�
�PON��4.q-�b���������'YR�^Ug��+��� �4���e'O{Y8j��#x��Ȣ._6?���AMb,�),����&IM���"#��c".�m�3-7m��~�_��Ɉ(MZ��n� Ez���2�)��$�f|��=obhӠ)I�݌�o���ޚy�/���D"'$��c��`QR�|����$t�	���.Yӡ�D\�����DYo_���H����s6lZ	�::&c���8��3�h��W��+���X7���o�/���&&7(�ݹ��{b�.k{ʨP���%é�)X	(�
S��.͆���G
E ��`,�R�,��5S�kN� <#�=���cP�*N�e��zFP�2��U��ٝ�^�k(��L��;\:RU$���cE 6���
SOat���ք�X馴����
�r��68՜@��ͭ��<����Q�K��ɠf��.�[��-�@z%C����kWm��xU!��d�^�喑L���#ƣ�Y��
t#Ǯ"��e��Z�H��F%$�*Ã�eZ��d����T>��IB�ǫV�5ǆ�H�L�=G��|2�]_�O�'jZSI���C�i&�1��W���q��y!ɎM����P	�Q�^
��*:b�&F�F~
��A@c� R�������3��+F.��U��V��&i{TO��G03��*Ȧ�'�%5�i��̦:1�1�D\C<fAO��/�������b�m�k�B�B��#Ĺx"��X���D
l4�O.�(T�8D���(�$���&u��ٚͿ�������:���x�ð�__�ۍ��Qc��*��\��%R�	5j�� ���3�	ѐ����(��?��;Z��\~v�=����Ir�� ��C���Q���X)��WQQ.�t��R�	%�ד��>g�.��|>�ý�[�����Y+�Sf���{��y�B�0��b3�$&�^�JHE,���TA�9�l�N7`�h�&�Ɋ�㞋���B�w%�]��C�hM�L���{1BM#]���4��@z��$,�Ì�얇�T)�Q��ap�GG8}SR��ɂ���Ő�*�T��'�J1�`�A�><LD:��|x!d\3�Q�� ?�
ɅZX��D%^��+_ a�^0$ �Y������ߦ��0ch��])^��q6�9U���ni��g�µ1�dS�ĘS��,�������@���4��~u���������������'�?�LhFe�����T��ƞ];�p�5WK��h��������DKL�gv��%�;o��	�|3;ϯ܎�(x����kC-z��J#|Z��yD���'���{�2ޢ9�ĵz 	�6U�Y�)�l����7b!�MX�G������C���;򜄮f��LU���� Kc1������*]����OZI�U8���"�Ia��(�m��(ds0T��S/0
<$������Q��5|vنB�9V"�Q	�{s5�Tp�lh�`�MG8�1�.�뗒�z�h-�S�(i��h�8q*��+7�4��J@6;�kA���t3��a(�S<�]!�����!w�
`�#�i�&;�R>�oH%�:'Fg�U���бY	vv	��ȵ�KC�dR�!�gK��/"P� ����i�ȅZv�,:��H�S���0LN�1آ��l�E�P��gWON�� 07�
�bZ���i�DtK,���Ɔ��%�� ��j�.(�)xyQ��;����(����X��,ƴ�
�k�Bd��L�#�(hiLC��سzԀ��A��Ʀ4�JY�8����GL�����{���>.��W
��Z-u�?��x���htߩ~XХ��Ǆ"� ݂X;�f����^��UCٌ�a��$a��T)������*��!��8I_KX�>��>��r_�a��5N~��r��_�\C��k��Hp�$,Z�B#�����f �������*�&(������k���u���H!ڄ��]�U���B��tq��&<�\#�chR�I�:T���iP��W�����r#���[ߏ��F�;<Q��<b\R���"���n����*f{@�0�kD:���e/XHx
c>yH2h$$���_�}��Oq�����}l��Qa������m�����[�s�c��8b�$�w���
�t�C���Kz�����UW!ޘ�K�Ų%<�v'�3B���C'��G�[�n�Qǟ�I�g��7`[i�x3��
�i��I�A��@)��s����i��2���~ņ�<���3C�5�@7�:az,h����y$�C4�d��u	��2(�F���wr�R����eDTDj&
ݛq�!�q�Qsеe;x�1�M?� ��ޅ����}����Byx �G'��O-�ޞ^l�>���Aנ���6����UK��<�Q��,@�|+�h$�Ш��א�n�$DĥM�n��4���
}�����N�%2ºW)uU"(�14�d������(�U�\i>��Z*�\�Y X��+*�+�<b�4KL���5����&��9!j&[;�sT]��\(N�[��Q�1:=2��*�d,�����`54�?�h�BKa�gb���zC"���AQ��j\M�!'l>��#�Gh]�
U^K*�F���{�4X�ҧ�+��cgfT-���6��0T����y\`���h���@GKB�"��k%t&+(��G�5��jp-ј���_�P�4���`V�a�2B��L�FUS�C�Y3��A����h�mőu��)�5��Ƚ��s>.��W
���Z���o~`�7*k��\���՜@�C�PΣq����b�sk2��*20��]�+^�_s�
B8��S�H�"���5�����ˮ�Iv$l']"�܈0|=�m)y ����a^^l����B��	�=����(]�Մ%IhP���Z�tn�����>��x	���()�<�C9g��1G9䥠#e021�ر;�)PI����F'l6�7 b1	�_zq��$��dn��9y�l��M���"������N(RF� ~/�ȒVReZ�$�ߩ����p�Tف�=_3��47a_���02����/����1+>Nå��v����w᳟8�ޭxk����u��v�Z�[w��j���6
���(�R����2{׼��~'�y��v,�Ћ��X8�����Y�%N�
b��P�V�#��Ʉ�W��H���ԅB��')e��w�����A��VQ�=TY�U���V��k��̼6$G�p,�����
����pwj�C�6�A��#B��r�Ӎ���eЙ�K�>U����Ȗ�=�МjEa8xy�e�u��?�D,[����~(�CQkhC�FK*���� ��~�y��ؿ��'O���X"i|G̙.FPTL���p��/�@5�G^�-�&|C�;Y4 �+/:kV���/�ęg��'�I��Ҋ�سo/>u�qb)��w/���-M8q�B,��^\��/b�@74��y���s��4^x�e�z�Qx����ih�A��_��w|����	c�f����
�jJ8�CϬ1&���N���<���X��
���O�}ܮ    IDATa�As�St��O�
��UC*�=7I�lv9���s���<�3�ἳN�-���M; ��;�/�f�)���=�B�t�'1v�d�����b�_���H�u�����V,~�ET���U��8�_���h� ,z
�z�]�}�'q���E���xc��埠4NF�~�A����� �B���o��s�>����1
��_s��♘>�@����m�&��ꋰwh7?�&P~��8�������k�_���������Q������,����_)�;k5�W��mz����Z����s�dA�m�t	�z>"*wr&�.qc�bux���3�:M���ek��y�k&�dC7cЉW��V��e�ģ�}8�H5��r�-]��b���hUAM�=&D8�ք�[5(zV:i�I�ԵH�@&�V��	�r�b��?��
����X�>1�Z���8�u�<C%��+��e��ɩ�6�|��bYp9E������h$S���e�Uo�z]�U�$E�� �49R��7s��ڐ��lA�QH���H�>٫��'$nd3���W$��&���иgg�g�p)G�V�0���A�E�ʈ;]��:&5(����k�j�۰F:��B'��	q������7��h��t�,d=-�I���8l���D:�v�� ��K	[�t< (�^+
D�C7�!��r��Zp¬�UW]�9�O��
�Id��F��0�w��P�6W�U�C��ahR������HQw5,��>�)����u��cf�W?\�$��&$ǖ	Sp��oC�7���`��ڄ��-�Q���LK'JH�����*p�p�5*x���e�N�ͽ��Exb�;X��P��?����`����B�j�#���O}K�w㧿~���pi5j ���p՗�ƥ�����w��o�os�j���p��Yx��p�qs�q�v�`^^օ�������?�c,^r3��T�O>�k��R`��`o�~��ۧ⍷ע�g G~�{�y��'���m8`�d�z���Ոd:��U)�!���[�\�7�@Ͼ��ف���O.�C5ւ�,~�yF2!��c�/��<J���a5�F�z�J	J~�x���ƅ���g�cҤihJ���g��[o���7�,݋�~���ߠX��3F��|����e�V����;rxd������l���QE*(�ٝ�慧#e�=�,��g-»��@۸�@��n���5�@ʲѦ����S��P	��o���kp�9g���mX�b�ޚ��/��g�X�����U���kX��l��go[1,l���k�Ŷ�Z:U\��7��]�f�:�1���~\����Z�f\�x�����S��Q���$C.�j}�8 }��J�"�	��8m�E+�*,���z2q22U `/$�0��F�wz�6��V��$@O�d*�Y���������������N�L��"3��� M2���f��ɉL+H
z��\��4Z%l+TzZ��8C���ߵ�'ta�K(T��CËz!�W%䃨Ӝ������ܣ�	c*�U�%[ bPݠ3Z�ժ�]8��������b��,8���?���dE��0X7L�M��iI��,PmDja��C}9=�ke(�AS-8�\2ݙ_����Ъ��/\���珰��T���@څ��dp؄�>���>w��;�EC�h�ܹ�un��W�������A,~�t�?
�9���T���(�hR�BU����ȨB�����Z�Ƽ&J,�x�'ǂN��d*�	j��C����zY&tS�?�B�Q~-����%R�id$�=D�]z��-(�.J)��6��uȄ�gQ�����ϗ��d�طn5n��E��ٝ�lj����>4N���wߋ��et4�A�Q��㖛�ǢS�C����҄ҿ����A���nT���@v��X�"^v�J���W��m��_�=�]t4�x���P�2.<��}j�/Y��Y/Ҍ���R}h�����oal�͍q\|���88o�(���38��s���Wp։���~�8�"��:	k׿��?�:�x����b� �r�Ex�O��A��aG_��N;7^}���]]�r-���#N�7��O��}�+o�,OKOAU����O�v>~��Gp���~����q�G���ߌׂ�>Y6��^&~��/�'y�W���a_��'�� _K"jX�wo×N���}}���xW��M7^�?�}
�a�E7�t+n��F���sx������������㏃i(غo���=���&�����!�Pڷ�^�|`�=�����O���)@_�����F����M �8P��0����[~��]E\u�M�0il#�v�W��㟯��I�-�O�v*��"����?�/�sz�9|��;��G=����/��E�X�� .��#0�N�0w�5�3��~xb�|��|�r�77�[KV�{`�3s�"��Cͦ�8}�HR�"�"$� _�a0F��pY(�K�J�D�lY|�I
�G����e4�JX���]���C���P� �,52B	S�6�DTj,�FO�ߴ���N֮Ii�L�U���Ĝvf�!z�	a4]�T�\E��$����4Q������Z��	�Ӛ��������G�O�g�L�#lx٭��p`W����Ua�FM2�=ѣsP��j�ə�"k�����׍5Fvٲﭿw) "ocQ�O�R�HcWjN��]�����N����˪Aԩ͖FɃf0���Ы�&�qIJ+`ښ��E��j�m_�'��Ǒֈ4����K��{��3f6��iǞ�_��V��%�Vl��koG�c�j��jء�.Պç���?Ӂb�j�?��	�h�V�|�QCd,�B�cAg3(��C�b7`���z�ՇJ��&���I`t���JHTa���<%a�W�v䞑����5�/KX�Q��(�aT�v�?�*>sj��� �B��q�y���O_�Y����<���8��3q�QG!�zH�fP�S��{��=o��4y��X�+��6څ*a�����?��|;L��TL�}���]���F�`��V�����?_Z�X�XD�1���aB"�{n��#���o[�sf����ϫ�V����~y���U8�3���k7��Ϟ>}���{�²u}�������~�c����G]��O8�_}&6�[�y�BwO={�I:ܭ��n��v���0n���7�@����<����p�}/"O�?�:&�k�7t+�;��4�x
e!��P��������t��U|��?í�D������K/<O>��>�v�`Æu��g΀e�bl��_܉SO9��wc��w�o]�>�-Z�V�Ě�=xcs��jb��[:�ۏ6���]�L�h₳/�׿�i�p�BrYL>��r��_�j�T��
;�bN���~�l����ށ2"�=c~�����/�/7^��4/-�V^�?�<z�ϰ��?]�
j��
�v���7_��Z�?��Nr�����������}��jf�ח�Ϳ-{��;�9ñѨ�>B�5GdX,�b�@�T-dtr����N	au��0�@���i-s������qϋ�Y�J8)��,B�Y�`Ҵ~T8��d3y�Td���i�-��N)I5���TAѭp8����4��3��
��_=�UQ%�ʰě9�
Pqʨ�V�0CI�[L��>"l>��e��p�,3؇NU!I�CX�e�#�Z��--LJ�l�B���,��L*S樑g�`2Yp�Pv��;�x0�5�!���KE42�ɵ�I`zR�X��Ưר��44T�
�l�x=h.B�_��o���c4Y�ټ�6�tc�r��:�@���(ܫS�G�+�A�&B&PP��1���c���W�7���W�;w�DӘV��Č��_�&Lj�n�K�_?9#%��T���H^���+0kbGZ�V�kc��#)T��$TTͳB�� ��N
4:�p�5�(g�/JaAW)�e�Z*�f-��a9�p�T%7��)�^��s"d�$b�gh���ū[$��N��k�)���ұ�8�j�~�������ƞu�1y�8��.���`)t��[�
;wm�M��>d6��F����c��͸���A�L@5ƴ�]x��b\ܗ��Œ���o��G�!Sp�__G����7~����E��6������ᩧ�Ǻ��/�?����ҩӱ��������K+7#��$�+^[��9�<�,>wޙh� �e౧�Żｍ�_�4����.���c�H���x������C����~�s�4&���'q�eg2�C6p����;q���ż��<�?Ĝ���.�a3bB+}f� Z�w��ۂ�qQ��o<����!5���z.��T���T\��l	��o;~x�����9�|�����N�c��1�?��.��<���N�Qَ̟�����`�;���+������U%\q�0F͐3�t�f�q����Cg�����f�:̙7�g	�p��A���"h�j��W´����Ɉ�|JI#<���!�[�:���E���Zܿ�
���{vn��.8?��^|��b�(E�.߸�?�Ԕ��7��{z��z�8�kev�45�^���!����~����%�����CX����HAg��*2m)�`ܦE�RD$C������P$j�yx��!T�<��
j<��Nβw��^��Q'�H��$�VS��%�ĨV��@B<5ɺ'z�T�.�48Ur��Z���j<:X(�"E]1%Z51�ʁ@q~0JД������#+W�pw����#y�u���b9�P����y(QB�t�2�D���CcJMdhۑ�_{���W(��X��8�YV�A�g�L�
߷����m-mm�S��ݥ)� L�"h��˓XP�֜l���x�BQ��#�+1UD����X_���3�M������Ȃ�B14�����2�sp��6s���O!�;���ZXQ{X�e�jF����~{
Q 9F�M&JP>��-+m"&5y�lp�B��\`��.ˀbV���O"u�t$�!R
>C4�1�W��R
.�M�l� z�^ぼVj�}rE�
8:B`aw�������`
�&N�5��ڋˑ|��W�kМ
��Ø7�s�Ű�e
�M��D�¾�ؿ��d��x���	0q�,<�䋘{��7c���I�Nd*Ԡ�+��)sF����*�ĒX�j5�8f!��ن�q��y�v�܎/����x���w����՝�q�N��T���p�a0�a����q�'NG�=��� *>�~�z|�Ӱ�՘8��-��a�6,}m�4<��?��_���V�ٷ_�y睂1���܊h��o`�1���ӏ`��ÐLe������E�c������b�&Z7��:Ŝ��6«hQ�8��lhãO<�={z0s��y�<l�مǖm2��1Q�MQ�H&����X3�8l�Lă*���8drS't��e+�6����e���4,}eN8�0�ūb�iػg?^~�E���܃f
oh��M}xoKԦIp��� 2�m��M~��aݖm�y�<���q��`���6�l-��>b�q�I��y��?P�(�`�045���LÎ;����Î<�6�B_�6�r�X��*�Iw�%���{�+yX�9�@ӱ���س{D2��t
8�5����Ŷ���c���܍�>����m-Aȝz�Bƺ[_�W�NM:��1��Y�T��P�M�kܡ���a_2�9�q'/�da]sҭC�r����B�T�+�YJ�|�0�C�M��o�ot�2	Dk��o���h0�Ͱ��z�s2�8z��9_��4�A�C�b#�0����a�d���&Ҳ�%��L�lx�g�qD^g�"{��N��Ub�Im<�%11̨�	��Wa&"���rn���Q8CEDu)˂TD�J�7�u�@�FyNņ�ޗf�&�(�|���J*�s�hT,\	�ۥ��)U�QFkDŜImH*�b���à�@��A"݊J�����0��!��&Dg�Q]�2�������8Ї���gQ�{�!2��P����҈�"���hK�@����É��UV24��|O�X��s�N�dl;�:s�T{L��])'-�;��G;����j�.��Q���狢�`�b�"a�@<��*�bqh��JņG��Tާ�jDx�}y>(\���0ΓBh���Ϡ �������B�w �x
�ᢥ��J��Nٌ�"o����!�Є�ֆ��-�!�̼�B�)@u�P36�J��>����R^Z����X&E��PbX�d�@�Z��B�sPR�oI�DQUE�D�B	j����B�m��\6o��{	�I�W�2�E��=+&R2/?���(�Z#LӫT<�h�oB��	n^
99�D�!�*�ǅ�E`%҈E5��0k�Dg��I�e���G�(�j$�RK�<��J6"V�[���x9Y㙱&����a9�4 ������F�P)�yԐi��p�c���zO%�He%� e��ȁ_D��C`��kH�9ɱ���|��R��(�	$�_c��_���]/"���p�k������YB�V22e����`Q���H�S`���^�	=C)P�qdk4��U�h�(sL>j/��z����������8)��� g��7�y�	�ż��#�Hbحam_�9,4H��H�'R�U%S�,dj)���5���;�����S�>��~�&�F�BZfv!/�dNz�ړ:���uNĠ�c���@C+|-q1�UX玔<3�#��E���0c�X���Q����::P�IJ�8���0��nzC(�5�NX�򇶖$�jg����b1vnNa �1��8'�Z�B������2}���e�*�����DC����WC4ӊ|%@$��O/m8����%{��z�#Z���2��lZ��̞c�L��3�ڄ��2Ԙ%9ޔ��fH�ߚi0��� Ԩc`).��^ă2ہL4&���ף�F�Fǡd{ho��o�.$��P5xQ.mG�*�x)ņ�80�,H�@M��<�F٭�j7@!$��a�y�:IO542l�.JͶ� =�?4�\M�מ9������,�<��ە�CA����Bқd����䄐_2�C����,l�t"&�#�E�eᣅ����$ߣT�1d�d�e1(����J9R�duE�r�b���`h)р{5V
��-tw�4���	\��@��V����h5�I�P,�E��?�-�ڔDvp �L��p��h"�R�ī�L�k�Q�
t�X&�f��R�Ascl�����%i�c�$t�BNe�H�&�t<����6�
|���AG{#��´2�9P@9�P��?�CÖ���)tT����W�Z����"~���Z�1$��� ����.�4��[���L"64��T`�<'X�I�亱����Ë���U��L�Q*���#JF����%�0bPOn��ˢ%q��<[O���9!b�L#[�#� �l����ONQ\Vp�dM�4'"�%�C<��p��Uf"&)������bD����$�������s��g��CU��Kc�Gq�8��|��3�?J�����܍������7���F(�,�bcJ�8�H��ޠ� ����tr�"�����u{�����A!*�V�p{��3}�-IU�t(Ll�FC$�rDC-R����jF%��%]�X�8H*.�
��܄m+�����y��􋾉W6���\.�f�N#��b�#�O
�|0���TЖ���Z���E&�����Q���68���i!s9,�uz��F|�	��ؤ���]�]�l�d`��%������Hz]B� ��1Եje���@�4�Т�"�+nY�0]��D/�j���>	%G���%	3���l1=��G�t9�8�Cäh�8t*���^���L�3'�x���ؙK@���T
�����	]��q���Z��x�I�������aVg
c�*�v���ń��WmE^�?҈T�/�䠋4,� �x�[@�菜�$�W�:��èVU�n�8�iFU�1�tǢ��pQ*�$����N'�8UW��/�    IDAT�Cp؄1FR���	93b��v"L�L`��ʤ�d<��L� #n:�\�~�;w�� ��Ԥi�ǁN#���T�b��71�&bqN��J��ƦD�]~G�+"���r��\I$Pa؇�!�͢��)<�C>�"�p<!�1[=O�٘�Ze��y�G�����ѻ?��əhN��P� |'ݬ�H��v
D؈�9a*�<S��n�����P�80�(��fV܄R��+�D�1m�X�T�x9q����7!����S�@t�T�����OzLx�ɛ��$��2A;e"_��#SA�`�62	��~���Q-��)�+��c�1�+0E�~i���a1�*\��H�6b��XbǳE�t�t���0����B[ߢ�B�g����j�Pѣ밫
]��d�688�d,#9ӭ���PP�L5�l���JD�t��f���F�����p'���7��b���V�ZC�v��|�2`ő��s/\&**�*y��?}�9C����߽�+xk�_7�����?:��,� �E�cFe?��-`���k�[����]��)�0Fd[���ep�^��F
z8����0����/td'?���PsTDA��J�4�.�#���c����_�&^\��]eZC:<A�E��=���(j�����Z?�0���������|�2l��5.�V�8�����>��.;��(G~x�pr�i�C��m��CH�Z�&��Eip��nu�,:{�y��� �]�E�����M��!h���L��~!�izf,��ǜ��ۺ���/c�ę�"Pci�=��d��6�W�K۩ e�G΂���q�~�"~�����/�K�G���j��N�$�yr����4� �i����]��bLc��f�⽗���W�Č�3q��/����xg�/�3m�\*E�d�V��"T���I�}���B"�L�S4�rY���V
5��Y�|N�����2:��P�3�Gh���T.��ĂLn�m>��Z���R
S��O�ס��K8p�t����݂�0�Ӳb2���3X�\����$Lwy�8U��1�Mr#s쓩�D�r�'\Zf� 7;��^��&,-�W�Et���aH��(����X	h�������bsʤ��1e��k�p��^-�`b����D��bb����T("��#W�Ivs�gMG<�R)�P��hЪ��0���#O#m@oo/⩨X�g�1s���/ᑯa�N)�1�iزq=jՒ Tm1[֭ƨ�Vd�6�D3jVZ���4�wH#���=���},da%��0�1�q�����ǭb���{#���1����_]I]�04��a��]IH���$ah&�J&Sm��F�=���D�������v�lW�^qdL�hmM`��m�b�(-1TἌՁ\O���D"-Q���fi�d�UqђjF�@rv/��
\���ac��chj�����j(x1�V����$#�͇��j�\��R�Pi�S�����
r�V=�����aq����9���O����t��1��(�RF w�_F'y*�`��Nj���;nE��q�/���ׅu�ԭ�ڀ
/NܶT��H��o�ꔝ�O#Edᾑ�u�5�1��V'�uГ]�ԊNoT�=H�Y�s�xm{�.�ǝr6&~:�o;���@��,c�N=�\�� 7@ȿ�����6эc�Z�������/~�3X�q;^���8^4�b��|hZy�'t�d��`Y��d��Ϣ���~��
���{1wb{�����p����տ\w�m�2y�L����M�MQ�ߜDfGG�RE�H�q�X�k�yqq��0e�tl���5�� 3�`ow{�!l�=��r�v�Pl/�@M� 0-jb��1X��+h�0}j
�fၝL��n�<0���c�P@��U�w��KG��GJ�☹m�پK�y�g����'a���3ߌ��'�ǋ54�R��MW����1:G϶�H�#B���xJ%��|��	�mG��fH:��lң�
�'cZ���ɂν�AY����]h*� 	���׻��a�4�_��\!g�4���0a�LQ������u�^�ԥa A������@]�Ic���M#���s�{�h^M���98�ضe+��lQ!��"�ۚ��u�l�%��vNb��!�l�����(�rhj� �I�=�_�TC�׮"�j�]31�@�x���&�1̅WEu���ASD���؀cl� )-���"�H�ш��fs���CSS��
O�'{scF&�����1�Z�턱S1���}��0a,*�OqdZ�� �a£7�i��w@�;���F���jlBw�~X��b�%��>��?�hyJ�x��0U�b��(z� 7�(J�,L����[E2� �?7�#�S����M�i�Fܨ��K2��3Ր���"В
��$�hll������s������SA:��g�2\^L2�(�n�M�^�4C
j_��9Ñbc�BI��%86_��H�k�������:�m���Xt��H-����$������3CF�G���;�s3�x�e�R>�Nq�r��|�p�J[tZWF+�8bl)�hZÛ{r�k�3���5qa%�%��A��@�!:a�����!�|�C�аE�f�OH�s �:��U�A3}(n/ҵ>2},TZ�jQl��]T���p� Q�'R�N��.`�)H?!��B�d���-LmJ�?>��L����x~��01�����]FX�啇���>���k��k���D@-�ePEi�r�e�3X��+8��h����q��¸�ӱn�f,��C�<e�]&�TC6n؊k7`���#�x`yH��ؾy"��5���9�l��v5��+��4ȶ��ǟ�1��&�j�}�&����&s̨��g���1`ʸzsl�P5�� ���Á���#�,�h����E�C�jD���X-�ٝ1�ooǓO��ӧc��V����.�QKw�L~���@�QƜ�!���kͻ�̤��as�!�$�Q��bP
�l/��%_�ќs�p����Ï���p1$���@��-s���5j���L��|%�r$HЃ*�9�tKKv�ًɓ'íV���'������|���-�R��=����V�h�,��8eq
4�II�3�(µKhn�õ+p��.qW�L�P.Rm� N"�eJ������x2p�"�_E�\"U*�(�1�k�&�Zvd�C�P.B�+�Պ��,t¶��\�!#R�c�����S�s���eX0��9Nx7Aa�VԔ ��$�r9AZ��4�H]{��������dQ	�B�KGQ*U
�46��/�s��E�);r�ٔ�96b�$�t*^Y�16Tʾ$����QR�W��&�s}HF��!���n���`�g�pX�X���rbx�b��3�/�c"���KDo��!M�A�0ј��.`߾�hی� �݈�T`���D$.�����H!F*�D9_@kK;��rR�ӌc�|>O���s�T��ފ)G��Ʃ'��eaqكSf;��d��C��X����	xnj�%�ǜ{`�Y��7�������jv��X�dk��!�Y�F>5�eE�No0�THT�R��o�(V}�+:)��h��Ƚ:�'�i%��2�ꚰE�|Y�Y�oC������!<���Ŋ�~����b\S�8'KX�3����T|�����b�@�Le3�X�ʴ#��3:J�Um�0��^R�2��� M8��2W������	8�	+��>�B��o{����(tj������tIt�=�M&5�5D)�*�1gbZ�����q-bZQ��%�+�9�X<g}�q4{:j`���\1@WW�4I'�|2�z��؈���`��R���3劍�����Y!�`A����F�9H�����w�&{��8��L="{=2�!��%G) ���`�"S��/$L�c祥$ϧ4Q����ˡ=�cʄ6Dc4��b��^��+a����b��r� �mL2���Tv����݈)-X��={`5�`��V���IS���'�@�se�Й�-D�1�����,��N�����{�b��شi֮_/�6�/��<�Y=<�Ŕ)S0o��F/e���X�p!֮Y�GL�&�{����S⩧�����ܹC��ѫ��_p�yg�z��t˥�L��T��d�QGa��q�:�w��|2�A&ӄ;waמ݈�Q!��NY���/Zt"�!Mr�P�m�׏<�H��t)�U��>�T�IT�,Xpz�w	��T	��8x�<��z�46l�{�XDR�9�݁9��捛�a� ���b�	شy3�$��|X�)�1O�x�iS@ss3zP,AN�-��;O=���K~��Dpf�����i�1�$�'Kʽ���7V��^x�%�4f�����8�wdr���0�s��}d��1<<,AA^{��3ENW���x�+e|���ށV�' 9ol�z8V�^���0�V<L��z^��Zfbg'F���W3/�(���y'�p*�/MЍ�1p��2W�(��2�O:￿����i����9q���e����]�u�Y�~�%���o�V�ޏ j$$v�{uQVH]���?徔���W��X)�F�[������\��Ƚ��RA���-`kea�l�jS�A�hp	�)�8�gKR�n�+c�����b"Ü�ZU�xT�s�\��e#�U`�j�ѡ�R���.�(	l4Aљ��A�9���)�p2�kԇ1�$u�TƃF�Q�� �D["��D�B�qMtՔ5ib-K��X	N�hm� ����J55)����ɴ ��|cr$���;;��4#���g9$k�H���[�����ه�Hsf�C�<��0q�x�~�����	�-D4�Ԩ!��m;va�o����'ˍ�7��f8L��7�P9X��xg�u��l�܅�|�^�Ƹ���%�B��b�����&��È�0���D��H�*P��`Q�E�Q�DT�Ȩ5���%٭6���ř�0TjqxfR�Ic��RŌ��=/`���ud:�2E��&L���}}ؼi+Ra����B����W��U>�@2aa֌�8q�L�<X]2���+mٲE��2]F-�dKv	�]w��;M�n���l��޺u�%1���#�ݸ
��jkƼy#��\���{�J6�g�4z8r}去���E0o�\���"'ZEϾn�(V���==�C�?��,q���t
�&MBgg�y��ù!̜9�?�O�ڽ�xB>;l2�8���itv��̙ʎ�E�u�R$�;:��#� �+"�	B�F�χ�k�Y&�>j�����΁�Ax~��mx���;���L��e��r�����͛'�_V"���r8Q:^~u�X�،���s�w�D�ǡ���S�J��L��o�~$�DS<��GD%���$S��ЀH��܀c�>��D �������T�����W_�隤L�(a�*���uT��ޖ�fy&�\4557�>�o��R�.�ߡ�a�;
{������`��7}��tS�ѣ��������[�ҩ4J�p�C��P6�#�ŉ'%?w�w�\c�"�p�=��뫘vĩ��xc[�xZ$�O��KȌFJr`Ѯ�� �T��TL�h%�1@���n	�6���=#;����������������#�р�����rB�5���b��9�e��ǐq����1�S+�Yˢ#���V����b����Ĩt
���0�%��N�,?����B�sI6cx
-X�!�C�;��
w��|3�T���&��	����j���#J�N�'�D=t"!��[ŕW��hh��8�e�GX�w�#�b5�Oy=�\Ӽ�xN~����0�3
�t͊���������/}����/��>1�xy�r<��R����}H'(g1�JR��F�~L�>S��֬Y�
3�QÁs�g��wV��+�w���ܽ�Z��WoÖ�����`X��P3`��D&*B�4硜Ml�x�q"�P?--t�!2#�kf]��	N���(:�\|1*2�d����6�;���+�<v��cb�d�Di�|��*�ni��.���{zaŢ(�K�>s�Dc^{��ИiƬ�b��_ݫ��+W�-Q���B����d�?8�O<�>����=��mؼu:ǎ�/~y����wp��J��/�9��N8�����{�Q����p���?�)V�\){q�D"��`����'M���>@&��"�z�Z\���bѢ�u�V���f���d<.�=��)S�㎻���.���y���Z��K�K1��̯�sGT��p�����w���V�SNR_oO7.��Rv�|Y�ݳ[�>�$׫����i�G?�{v��3g��6���j�{��x��7����H	�f�h�4���K�*M�!��U+�F1��}�݇O8/����Ɠ�v��z�:R����P_y�����4���2ڛ�p�o~-����'E��?^g���ˁ�g#��ɽ ��H��O�6���a}���Ao�~��D$X8�¸��g^r�%ro��y}�
̝;��r��ݯ��\^'w���|��7u�t�V7\#F���;�b���1~�8�=x��ｳR �f�[ۥY�����z�u7�c���8d�\|��_Ƙ�Q҈�޹;/����Ow�?���S���T}̞s(�������CU�$��@,��͵'Wcaǎ*�����(�����zS��µg�{�#����onǥK����wA�l�HA��6eb��(B�j��!���'�@�G�����;rJw|����Y��VN�&lz��uܧZ�`� � �'O����
5(�^�aq��S�`�U��A(G!Ú)h����&��.�kO� �<��`�F!�)�4z�$Qz�В�hu�~���A�	PJ�w�!�K���q�CX>����ěQ7L�0�SUaD��aAW|D�U���0w�8|�#1>Z��UKq�1GaB[��j�����y��u�nܻ�A�r�'@��O?��>Bvr�oƂG������qЬ���k�@�dRϚ5�>O?����L?7mǶm�h�<�Jn�s1
Z�X��2j��uΘ��;����$�Y�jL�?��;P�B����	��d0�D܆.~dQ�.M�Z+�$�p���x	'=�)!�s����a|�;���W�|1�^x���
����fb�����;��W�-��'��X<)�Ҫ��y�̙-��T:!;DBۼ�l�Ə��Uﾋg�};w��؎qX�a=����J�����k�*�bف{&L�����G�Z��G�X.a���R4��n�K����&3l�	��U����7�y��*o��f}�-��W���juUX�d�sjoii��k�~�g������'A����n�A���E��������=��眏1�:�e�V���&�N��[~q�S~=��K�6����NiX���044��frvJQ�������|}}=�g�ԑ����mt��p����<��6�׭�F��{�y�R*�ԐN���k�knjn���\}�5����)�$�c�>
]t�4i��gҐ�ac�k�յY�W�;^
/�̓��4���~_A2����&���}�Xi��r����>̛`���Kb�]�9��_,U��ilj�?x�>���gE)CD�3?��}�(��E��"/���~�1<��sr���%��������>�h��#Q��d3�{�<���86��Ihj퀓���xd�fhVe:����K<�$�B�<h �cpbwM��"�2.۰�+8�%>�ϟ���HU�e�����}��zxWu^>�*���WA�a-0�O| �h��
h��E6'����q�o�YĬ� ���^�z��wı8��+��?�J-��x=o>�L� C�Q����"i;�L�❮2�}�B��;S�H�X�"�8
�{omw]�}_�=�g�)9�C��FA@@q`�Y�}Z}j�Vmkkm����c}k�V�*}lk��ւ� (�$!aH ��y8'g��_?�w��V�;]��+�}�������ắ+'T�������Q�����_�G-1v�laʄI:���9�&\    IDAT]i�Qj�E�g�Di<���Ugs��n�c�zϐ���j:�	 =�3�w������KG�OƔ��)\<�e���G�5u��}K�{����&}�˷鼋�Q74C<�|~��R1�;�,v���2�}�Y����_o����t�i�Ie56��D%�p�
i`���?��a̓��"��D�6];?m��QMuL�b!��,&L۵2�uf�i�4���X锅!�x���6늶JJ7T�|Q����C=2��z����7tՕW�i׋�� I������/h��M����+V����c�oFt���=�?�����J���ON(�ibjJ�\N���������f�&\b�ջ���Z�a �e�V�y�Y����ﴯ�_�ك�>�A��n���h��5���/��r�q�X���zO ���cco!]v��V^��J�y�{t�m_������Λ���ZCo��MLLiϾ��7H��a��~��DhW �qx&ac�����8��٫�K��ʫ��e�>q���,}{�K��������{n�e���?�������S���c�~ʽ�P8�#G���|����Y��@��������W~�s��#Gtt�~����[nQ�
��h����>��z���g딝cΙ�8t@>��ب����Y�N�C���g>����-f�ĺGpO��:p�:�C>���[�Ħ�l�s��Ώ���� ?�=�s��Dc�>I&�ۿ��n��v�߿�9G�l��[��g�{�y���2���d�>�����_��6m:���ѱ�:����h#�-��*Ň-Hg��S��g.��������,'38w�6���;C�/]���oy�O�3�K��׾��g�D���C�6�+�J�Lu�41$C��e�_�M�h'���h"10;ɠۘ�tmT�I{v4/��-=u�w���gu���6^{��柾�v(�3�-ԋ?����Yժ5ʂKfJK���va�>�v�(m~�ͧ�S<�V2�W{�HTo��J���D(��^�n�^~��;>��s��Kt�Шr<���zj2���!���r�Ⱦ�0CAKŹ�;�ts@�.��#+� �<���[�P�^S}�������~�]����Ӗ)4��/���ݴ�X���{�V�Y�����ׯ�c�=x�#����`���ٳG�Ã���X�����<�>���R&�����j���z��c�-?C��Ū������	��&&�Ne����UG¡��ug4�1��Ҍ8�R��X0��a����Q�í-M�I}����V�o�}��kj�Ұ������R�(+���ɯy�u�7�n�ވ�(�>�ȣ:t��'����Vn��_y�e�ˮ�r6� `�x�<�����\�g>��륗^p��m׻8oK�RN��a�|�}�_��#�MȶM�����,K�?�K��#n��/��d���0R�d��BO������� 2E"v,k׮�E]h�ɱn�p�x &��w��S	$ ��*ղV.?�J�����9�� �l��1�J��G}ԑ��ct46p>�9V�������q��@�bY=���F�XR_6g��h�kQ �h��5[u+�;�Bq˖��Q� �
S����K�`�|;~�E(6�&Xd�؏���'�4�"��Ȉ��g��QՒЁJ l�~<f<�ѱ1�w�}vY;.3��E���3�T�0cׇ����񌱞l߾c�ҁc#�Ӛ���h��nd��;�TAh��n���v��d�@��B_^S3����WX�dN���55��em�O�y���Ѳ��5�Rb��B�yii4NK�:�,#~�o�{�R8P]��U;���.Y�����<x���k%�_rE�������㱵 zP��Э�NY��q��܁��壳��R4�j�my�;ޕ鍨��r��V����U��ֺ3��S����1���-��g���S
Bu�2lu2fщ� 	5��T� P�st�;L?�F��tIO=]���?��k�r��^�]��|ޑ�{W �,Z�Aݟ˟��'>���Z=[]��_���̝��R�I��RX�d�c=0�1�C���RF/���Q�
U���Te�R�i��ߥ�F�ڵ�>��������_��Wu����ީۿ��w��e�:>vL�|�-�;w��Uk�آK�>=3���QMOM��-�ػg�~����t�+���}q��7_c��֟Y�ذ�aTm���*V���i���X��9g�]�ƣ0�=���4-j�Ѯv���ǚj7!@:�����r�l�*�Kfk���~S-3p�+\ڥ�m��j�vlݬ\�_�lV/ܭ|�O�j]�X�E���dYc	1v@�x��Z�f�� �K$��k*�L�#�r�-釒�Y*��` I��<%��۱����� 3F����3����`1<8d%�l_��p
�t���2�p���-���bN���\��8X�!ѱ?܏��Nv�s���x��'�p��xoÀ'�Z=����-�c���ڿ�r�z�wx`�Η����s����n܋�������f�gl�	�'�\0rf��k�@�KPA� �B��ew}U!�u�>>�`���r���< G�ţqhQ7N��[e"��R9 cz�ݑPX�B�ΑT�X�����\��sň��^-Y�m-�v����֛�/d�p? "^��vԏ)S��L:m@I��p�P��m�S�Z ����w����w>�{�xI��e�j�(S�t�Rb(�k4 �7D��M�ǻ�;=tL�j��D ��.I�����YN�����-��s����-{�a�w4]Fe$�hT�nX�:D��- �bX��)'{�T�Qu�td�E��c��͜�ֳ��J�-J��q~B/��B�1u����W�s��M4ԝr��F�K�G����yQ�P�~ٗ�|�.���{�h�t�y�ǵ�)�5#�x��
��.���������׾y��.�5�Ǔ<Ya�2+���&�u�n\+S9b����7N�D=&�8R��7 z���@�2������~U��Q��;���������O��V�^��rQ���w�b�j�^�Ҳ�Z�d��.�f�R���j �lgvfF�֭ђ�����/�w>�{��匉}�=?м�UH����xX�.S�Ʉ@ؔ�b���F��5uR��v$�Gk��4*$(���m��w*j�D;�]�)��J���Lq(sv�.�m7��&�S�3���5�_�Mo��Z���IRƻ�-֜o�1G���L�@M�-l&�1�X~�a���  �����\,Zp0�7���M�����pKÆ&`�Zۀ�6����-Ж-�c���L����X�Y��1�p�ܾ�~��fժ��s�~#ѥx:yZЀ0D6ӏf�<��5X��?�����d3�f&����e�R�x���>w���b��رQ�6�,��=�g!�b�w|��I;�����L��#U�VLnԘ�=� �v�cǜj���n�q��q�鴱ӧg	��v��n���3�����?`�/����vn	���)U�h�NuHT{��K���
���?f��ڟw�X��5�#}x�|��m��x?�����d�
zlydy=i�E�>uC�ݎN���8F �>� �#��*ص����]$�|�r}�#׷�ެx�ih����L����5���k�s��-��ߑ�����(ݩ�¡D��?�&{��k�qE��np��7��1/?�rU]������P����:�X�6�h"9.����-S���311h��ZJT�E4������%ƻ*�ۦM��:��gjǔ�c��F9	5*�E���H�5P*�̹����%,�Y��}��ϙ�r�<�ѱC������>�����W�������_b�?/?�����^�۷�4}�DF�v�zda��H]���bT䙕Eܤ>�c�c|�~wˢ�N��N�Lګv|L��Q�*GoL�9qTC鐆�bڲ�������6�;�E�kr긑�ұ�Y��e��5W�Zm�P���>g�u�^���~�!-Z�Tӓ3ꄓ�/W)2���Z�%M/�t�<�gM�s���+np1DJ�V:Vs�ٗv������h�@Dg�]����j-���f	�yk��ZU�q�&8�Ebƶ�_ߪv�hŔPQ����_����x�����l SC�-S��1�@k�řc�E��8=�f�$FQ�#��b��y�P{�$3�
��՗3�S�E�=�,�|FF8[��~)��� =@�O�3�VQ࢟ܝk {��Ϥ�v���py!� �@,���l\�<�Q$쉄XI�1�/�}�s'f�n��&8Mͮ�R>�bٕ�(85°3�+�*�mW�`��UAh{�'�$a��N���4DI��*EDk��=�Y���)�Ksw�����O�*@|皉��u�����3��U?\U�8:���&.�N�k��8�κ1WQ��F4�T6c���V�B�Y��U��YWٱgq�H܄Ld�X�g�B>����Xb.?n���2���}^�g������ܗ܏��QBG_�
 �GY�e-[v��x������u�AE�Pu<S�d&>���D<L�!P�d�Q�t�P9l)���)e�]0��џ_������W���ۍ~����ϋ�]�L[u�6@���@�!4C�SN妀@a�-�E[ű�d!	GT��e�J�f��������G{uꂌF_x\��1���UE���(�	�]X���D��ݪ�R;�*�HY���.��q��q�����M�a��Ĩ�+ �t,���h�ش��N=�E�����z��ݚ^��v��j��+X8�"�ߋ	a�� �Y�R���C��=�qd�F�y�ӻ
�ɤUݣ��--����%C�t�
��5}������\GG����j�����gͨnB 8f�ld.��ױ�c���OX:��m��Y���]����=?���szf�m}���6�J.\�B#�0�ט�tj���#>��6� ���k
P���p��|O_X������h�И.��-ʟ�^lA���|N�d��#mD�P+�-��h��T�S��	�ʯ�썫5�s1��?ݢ|.�F��z��Z	����Y��^X���<P��E�f���]�ʳ�c�Y����/>+b;'d�����8 �Z�^����N+۲�Q���g�f́�����r�Y/��'`���1ם�.��{���J:���}fL�q򻹷u(@YS�tO6	p8�<G��W���T*�a������J��k�l޶ۗw3���gW�(�I�@�J�~�vC�22Zd�d�5�Wo^��彀�kXV���qnL���׽^��y=�Q�I�F����ڨ�}H�Qn$ѫb�j���S}��Ú������H��9�k�FfN0���q�y����R����b �R�b�Kڕ�5dn��@���
�̔#D���Y�\I2����3*�]�K3Z�z����&m�yD������K���`�
)�,b	P<[��T�eS拉�R|��P� =ݭ낡x��?�������vc��շ4�k<�Id᭺#�a���S ;���Ex櫋�:�k��e��ʔg������� 7!�V���QSО�q�L��ڵ�ҭ�V/����W�t�X��"�*n0�`G���M�=�N��l��	s��ш�͆��陬[�R�TҢdj퐢�yV�:��ڹc��3�Z�j����F��QܹC�^>���(��U�2+�w��s�yn�.jO�SQr�6��^��(����T��pJ\�zG������n�Zo� �]�m�[/�P)�G���a���۾�Ozz�n�hr�迖l�>���&(A�k՚Stֹgj߾Wu�M7���-��,�e��gO*>�R/����Փæ��[�@���(hP�3#[XG�X���e]�e5E�q�rO�;Z����雟�4o����˴����{��7�h���L�J�0䱋`R��8�B7�f;�HkVK�ǔѨ�ܰB#��6�������U�w�@�^=@�3^f�ۗbYl1af��W�̧t�qM���3��,�����]��1���TEP�#a 1��f��m�s�zY��>��on�u������uD4� ��T*c�n2��@���={�C��w\� z�wXE�(n���w�p��޲��EK]����lˮ�pM۱ ĜS� 3k��^6�{Օrɂ��U����:�Ͼx2"ߋG�W7ˤ���9�Z毓Y����u�\H%�V��蠕��sz�>�4��W6�<������� 7�2���Hp�:.�U7��A�ީ#XPՉD���FO<�HZE���}���0;k����|�Qqu]����{֟�w������W����JbH�Xب>!S�D�)jDa�&:��c��hZd��51*�)%�u]4/Q��O��m����������j:�/aa�A�і���ݨ]��)S���gF� ;�����ۮО-�+Z�Qi��,��M^�b��pS�dLK�%�w�n�f��N�5 ���5JcJ��j�;
��:��n��ǒ��'�z��Zm=��sJe�&�	�Z��(6��dQ�������4Y�i��UnhH��9���x��;~L��yz߻ߡh��m/����MF�UPʤI퇒��ʜع!�� F��%��kG(����wjaEqlRT�򌺳���k^���v=q�����s�ب��i}�#���/:���lU*�������j����@X��h�����l8u���߯%˖��/|�V��wP��|Q����3_�z~��q�C�-X��Y�FLA-��h�������d`]��(��k%˅%K���MgR�J���׶��kn�u�:c��u׃/&�/P:S�<��K��HaH�F�`(�F+�ncJ�2Ǖ�t�e��J��P_6�p6dc��x�J_���/�r�X�Y<�q�ȣ��}Dg�~@<�ʳ�Y�- J&���7���9��p왔�{Ú��ղ����|I$H�ٹ����Yc{$4�?l���>od��;�1GX�(�@K�>)���ȍ�Fi�W1�}�?��l6�J�n�tH���� k�=3�xpK�0684d�>6ll����砥Q�B���d�%����\ ��=0��;玿���h��2b�>��
Χޗ݋�ٹ ��J"M�1�Z��ս}��B��6��L������mSl��Fv�����)W�s퇺��9�a��ƍgX��m[��r-�ɉi�"&���>�^�{*��R8�i�D�QĪ�	��m��GF�-o�A�د<7�b�� h�s�Bt�����x�ʹG�aֿD9s��Ͳ.Y�.���7����wt��]��;����Lx@A��n�ړ~m�g@�d�xZ��LI�TK����Y��������Ϩ������L�t�3���gu����r�t��Z�B3�����:z���{��ޟ|G�ʴ9 A�w\o�E��SF�YEZsĴ�y�o8r�cU�U�m�G��%���J�+T�Q�O�X��Z5�,R�Z��n*Ok�Q���:g!���PEi�����u���1t\��rE(T3�M�#
pw���[����qe�͎N�Y@t��N��֭�S6\��޽�w��b�G�e��b��U-EI�����_�Դ`�)*W�~鰂pZ�X�"霢��K)7���&�U__֒�J��N�O�X��ݺ.y��MG �8��#�h/�j�Ҹ�%4;zX�C5^�kמ	)ԧN@�w��v�L�:Y)t�p��4��f~M��a��|H�6������-�� "AX�Ips9�d���yg�Ǐw�P���R9ntͦ-� �/q��������Ik�7&��	���l�������Y��3B�Ij��o_�؝�i|.��|�V!#���T&�f�i1�g��h��ިW�"P(��f>#7з��+ߛO{o���X��G`��8��Q�� *آB��zV~o<1�Xܩ��&�X�L_*ͱ��~�i�DGf4|�e��d����1��$A�'�y��� '����g����C�����_\?2�h�r�r��F�4b ܔ��r=a��<�D6?�;�v�S�O���l�}w���,G��e��j    IDAT+��n۶͂6�ۙO����c��l/�}f;/���e�TV�Ym����Y��UF���Y�|�.��j=��q}{�Au���tm��������Q �9G�D���y��L�S	kFY#IŚe]�����?�Mݓ��5R�q9 Ž��<q�dr`66����9@�ck��6@w�ήH>�P�^�������������w��_����/ҏ�S�vG�Fi�)+T/�Φ�:ڏ�Kn�����|����������:j�c6f62<Ϭ ��Fպի5v�f���&�	�Pm*?�BK����-����M�Ս濬0���i�C�&r���zKc�(1�Тb�� �����PR��|���,A7.3Z�N�ƴ�zD"]eU�%͸��Tf�Ԫ�U�xT�zA�FY�Ҭ���;s�b�X$��)G&�D�a�Q��T*K��+���W�3��z2�Z21��lD����E;J�\�e����{�5Ռ�P�l�Q�p�J��h���	Ք6}���b	hV��3ى	�N��l��M�1�s�ÍD_��s`�G����V7��i��r���>�ł���"�����5���ղ֞b׆���lk��3@ə��)���V*s��8 &dj�/͵# `Q�����1�H�T"m�ۗ�	XX !�1�����+�3�C���ξ���=m����y���f��
��t�q�}�����Ք�={ݸ�������8�+� ���6���v���K�ιh9�A�h�ιf+#�^O4NC�:r,��fҭM7;N �s ݞ�.%�ևG[�������̹�4�L���7V�g� ��-��Rh�̿+#rn� �"`?x�����{*�h��t悯Tҵ�'@��ڰJX��d��
s�ѩ�q� [�^�_'x���1!;�}�3��8~��TN:���c�I�2�J���KV��ޫ�{g�׷oQz�z�I��Q*�ˎUT��@R�Z��	�9�F��V4S;��M�M�������� ��
g~�� �7����K�|!>���P@�d�|G�Mqd2�Y^N�����g��9�o~�w�;�]�_�������*�I�ڷW�ׯU�/�X�"��I=�����5�w����U4�U�0B4��Q�E3̍�Y��ȸr��͖w�2�v���ad)�S��5*������.�L��$}�.���������6E�isd#�Tf�Ʋ�IX�?B��	L��D�����!Ɓ����.� ���R"o�݌IնKY4���Z�м��:��J3��d�,�u��]|���KV�TL錞[��(��c۲�4:m%2Y3���r
"i�j
��
`�6��G��:��aG
�����Dú����s�*ڱoZ����J��uw,��7Mַ�v;��$�����V�~u�HV��NX�tƴ�±�ZU�"�������Z-�;�*k�`S�Us\����S�8%G
��C�<�	P����@ѕ�Y� -ߛ�_;?�������hS��J���5P�0��I
 �f2�$��Ŗ��^�/�Ą��;�]̠��wz���l!�Ɲ��L�@-e�l>���	%x��V�Zcr��A�A�yy#���܌֮Y�cǎ(P�8�;��GF���u��~�i��Ƿl� �ڷ�Ͳ�B���v��%K��9����XR�ס�ι�\"';>v�J̼�M���U�����fH���>zĀpg�M ;@Ŀ�?gY+����fBT��fן�
��>���0f�l���b�H��d�q�]{�8�- �����\��͹��H�W΁��ێ�@��=`�1��pp^	,)��xG?��wH�d����ǟ|����<���s/�7��۶���
�����n��P6��2.~����֞������¨������r5y��Ԍ��3�]���JG+�L���nH�tR�NU�DT�hR�FQo<e�t�'^#��w�s���/�1����7ۓ~m[O�-', Z���B��1.(q�4
Z�l��V�+��?��z�;����#�3zD+֬U>�����F�i#E�<�U�l�h��]q�jd�1\�:�6�
���v�U�JZ�z�Y��w@�T��M��"!Ma78�@��Vk��SEY�a���
wB���Q*?߈u̇l�a���0_�����Le�T�u'k`��\��t���ij*����r��X�4xx"�Wɬ�fbB��t4(��̴f��
�q�$2��M9��F��q��q��ɔMp���ꖭ���|�I甄�:|+���&�RG�Ҭ�����_��n=��۵n�2]~յ:R���V;�ge�p2�vu�ع�zW� �v��6��u#O�ф�M��[��M��$i�QS �R���}� ר2�R�[���	-�5oN�?Վ'�6�e�7� �4�!H��.���A�g��9_�6t��ʢL��>����4�e[Y�
Y��3�H����rc���~6��ї���[72GO�L0k�gX�,�.�n���|9�ZQ7�n�:m����{��a�.�����N���Z�4ϓ��{��Ts.��"���n��_v��޾�ZZ|~�Νv�9g�YvL��x� ;׭O>�7\�����7�p�2C��J�5�\�|���{���zU������}ᅗ�1��v9�C{^}�>����x�s���:㌳,!��ѐ��	��l6gAY����]o����Y1V���o����� �͍���1�����[������JgS��O�*V���1D���+��~,T���������c�����������*(ݮ6��;����{�ss��Wؿc���QP��:�j˦s��UW]��<���|nZ�H^�X��m������"�����M�qJWJaAݩ*H�T�&�fu�������d�N���J��j\��;�7����P�FZ��\�n�GF:V�iꝮ�є�S�Ń���ú����}��r�E��������L�_r�rɾ9�'�ɉ�ze�:u�j{��z�M*��j��Y`);%5S�X�����,4s����C��ʨ�E�*6�J�(5�D�䈦*Xb:B<����O�f�sG�L��D�)%�i�P17_PH%15Kh�G�>��'z�e$�x(�ϰ#nQ�.
E�T���z�T�3���B��*h!�T,j�n���w�3����i(��&
/X��'s�o�z�q*(8)Y���K7�L'���1$k:sM��.
������-��1�x���/Oi1��Aub�;���M�G�'�HסT[��&O�����4�j����ࢁ</{I��)>����k�^�3ڸ$�5#1e�gƴk�Nŉa�g���d���P���|O֗zY�|i���ʭѨ�����p�Y��LY0����ϒ1�1&�������e������|�ח�}flb)���F"�K��&7w�n��Q�6yos��1O$�0i�u�V��`���� E����:�}�27 0� vх监%�s�ݤG��F.Т�K���\�`�6l�`���?�k�Np��! :��M�d�G��ڹ��d˖-v�	>6oy�)�Q������5{ xb|ʪ �_��C�s��l��v��&m���զ	�YY��wQI�?�Q1n��6��u�>��=������z�Ǿw���M����4Gl�($3�t=MtX�<r����{�s��%-��P瘨dp?z'��;v���U�_������w`0oA"�~X��]w��z�;�Ȯ���=;��-t�HGx�X��M�D;a7��a�X�gX�ڊ5��`\�R#Q-�W�4�K��?���ϓn�N�h�]_�k�����D�_f>��g���Q�
��ѨHq�%�T�j�#�֦4���������]���_S��q����uӻޥx�E���(M�I���k���Z#��/^���k{��sx,�r��X"i�M��S�l�-�ʫ�訃0B(�����[��Z�H2k�v&�W��(Q�Y�k6�F�`�(fܧ+��U��W�[R�N�[v��S)J	g�j�\��^$Y}�&}�h��u�Y#����F�!e��X��Z��ߙ�N�c8C����
�0
h����;i�nǍ�x�:?"�[%������<&Ub
Q�UA����Z?����vM��iϡ��6T�$�˪Bxr$*xq0��Ȯ���hF� ��@����~�L\��֩T ��Sr�3�0�F� }e_M�ek������-iV\y�Lȏ#��x�S��<�{b�'VI��z�,�.��X��9���k��9�uzm&L5Z�9"��3b_%� nca�yx����ܽ\�/�d�O��e�^4�K�� ��-�͊s�b�`��8@�@�k�.ˊ��"����)����XDO=���9b>��{l��po{��t�]wY����x���[L#�`��( �+��j�t����?����8��q�F-[���d˖��ח��F�m�a��R}�Z ���Y��Ęm�N�Tӫ��m�O���2<��5.�u��v������|���y���z���+�)�J�N@�+��5{�U�S��3�|��ũθ5�׈J������<��p����l��\qU�.P�8�㣣�p�����h�Kc�Ǉ^V7�ت{|w��Qq�XG�R�!k)lv�X\co�zx�R6b��D��}��ǣ:+�����?O�:� �ݷ��؃��e(�
@7Õ�"ݘ:c/�jA�pI��I������
�e�����>�n�]~�)��T�-�ҕWcq�H8$��� �h�W��2�l_�-�L�)M�`eU"3=�񩢦''��f"i�=PX V-_�:�O骫���;�iɢ�������(^�cb`��md�B�#�DՌ��tx�*�a�&"
��ݦ�	P7�&%'�I���S���Li��pFh����c*���@�rG��#YEs���@���eM-�g:R̬h��ѵ'�M�t�R� ���|Yo�ܤ�ٽ��-Ņ�8�6��S�KX�<9Q��dG�FHA<�h�@�5
J���
�Ê��jB����Zn�Q(ém�Z�-Pq���ؔ�q0���9@_�����H��҉@=|�$�w�_Mv�}���"��ǎ��+��g� 4���:n��Dxz%�/^Lœ�~APs���I&���a ����~f�}#;���o �(8?N����O~��>���\y�s�=c !�j�rʵ|���^�{��Ƹ +��f{��;76��dӘ���s����~�3]p�E:p����)s�|?`C������aH�����Y��U�,������O�y���~���st��A#�Q~���t�g�𡣶O0���l�+7�߰V˖����vkt��}7��ι�}fλ'4r�9�~��s���|6�p�ܾI⚵������3�S����D��&;�|�b��l�o��r��^�������/���`�m y��<R9�x��ד���mL�:�T)�l��ʫoЖ�����U'��}D�J�UC0�#
���S �V{V+������{�Tu�eoг����;2���]�˃���tr �k��K��;���J/�O�)���y� 筤jZ�/�"%�I�,k���1�L����֣��UmZ3���x�=̏m~RW��-J�2e�W�a^��ў�_�ꕫ�/w�7[��?8�nbD�A���Z�p�2�wɣ�,��f�5;̻fT.�j����r��������a�:e�I�2�:zd�FFʕ���X�7]}�~��C��C��«ޫ;��k������O
�խ ��0�i}n܎j%��VA؂�=:�@(FѴ
�Jfbf4S����XT6PQ�ẑ�X��V�a^��������N�R<�z�@���gN��d���ӫ��K��yǢ�V}~D�]&m�/����T&�p�q<���_��	B� �nuժU]=Θ�uÐ�S�~#�A&�|�{�d鮂p"�G���0��s��2~� }듏jxp��y	�.k.��}t�ȃ��o��kz������،}/ 4 '�^M���~�r�	�8V�7;a�>�,�{<���a��Sj����x��3�������xg{ *�A��b�r-\8b�K&�(\x���w���ύ��%2;���fܓ�4<�=���I뒋/�}�"�x�ᇭ��6� �?u���Y{��4�e�s���p��}�y{�	l o�^�\۶=e\�{���Xy�9n��6��@�\��;�j �?��Ic�s�<!��#׉���':B����g�ݑ�0&r<����,�D� _ ���{�{r�^ԇ���q܀1�ʹ ������l-�Uj�������
�S��*h޼!����=	''�L�ޣ��U�ˣ���[��8�t�z�a�;n�2963ލM�E��u���e��o�3��o���o<S���41UֲHT_�������I�����K���c�E�>c�����aD����ZZ/��sOj��/�G�*���%���|Hw����yk���}�&���������|����@/f��+/i�)+���m���!2Z�l�����^}����CG�
"�0����j�DX��Ԧ���+_��NY�Z���ء}����cvv=�n+�#ǎj|��κ�L=�c�>���ԯ}�����czlϔj}*#;���F=�h,�t2�fuZ��)�S72�`�.�F�
@V8���]�as+ϒ�;Vv,1���I3���ˑt)���i:�e�˰���O��n�;��^�����'@�+�%��TW�V�I)ܜ9�pN4�0�Va�xoՈ��5ٶ�����tw>E���8�!t�;ue-�]빮�4���t�%@@\�]cF��'�qE�:�I��5m{�q�V����:E8������9��ۢg#D���{�9��wc76yOD�lp���@�(ZO��dNY�}i�Ϟ�~?KH�\��Iyq_z��$�E�˿~ޚ�y"���� �m�p%��Rt@�������N\���y��{�G����U�l2}J�7�@(�{��j�� �e����c�J�۩&�l�Hz%+�cM�9�ǹd�8���K�/��e#���}�Fy�}���1/8�>�9{�C`����/�)��	��g�}��+��yν���3Й��O�������7�g�U�iೖq.|����<@�d��3�����{���9O�c�P�9�x*������@��&��Vvj���~�O��dK��|� #%�6A`E��&K ڦ߁�E(�����xݙ���3��ۿ��r�ι�J��G4>YЅK��ӟ�1~*Y�I�������?����w��.�X��Sڥw�FH�v]�h]��Wd����+�ӂ�+��u���C/j��R_���>�!=�o���z������G���/�B!DW,�G:*��2;6����m��2b��˭����Y�r}�
��T�N��Ra�ƴ�j�A���V�_�\���g�Ñ�VӞ�׍o��J��3�[�ѣz�'5v�����`~��.;_��������.Y�` �B�h%wz��_�YQ\5-��?C�YU�@{�ul��*5�/�T�Ou��x��v\������2֦��	dV�-�[{Q)�l�b>���\6���[��R8$8�^N& v�����S�S���t��~�f���LR6{�"C���Z=w��]�W�-N<�i	H]nn�Um�S���D7�3�ܶ�s7�h�.,X��w�h���zJ5�Sz���V�Вg�����'�,ƞT�2��t����m}�XԲrcU��c��{<���	�L<I�m�C�����G�����#S�験Y�̟�eAgy����2u��	]F�C�7�����X�	4 T�1۲g�G~��)�y���Y(=x��;��7�f ��g�
(v�s֣��^�m�B>����~������M��VQ��1�O����ݔA�T����+�ql�5Y��iv|���ȞL|/܃��	`�l��l���s},���md�`���{�;��[&\w������	�r��Q|���� (�O�g��=����g=�^�fl|J##��fw��aMG�#�}�����q}o��j�a��J����f7p;�I��h��ZsB�����7���Uˌ�K    IDAT�8����z���KK���}�;⧞���D��/ߕ���9�]r"��y�A�^W$��O?E�][t�?|Yk֬�~���n����Ͷ��R��3�U�j�*�Je����:�|�߰�;䒎ʥ��g�/]j�M7�l�;�c�ϰZ�TarzF�n<K���*��%C����t��w<ܔ�-^�o��w����2zn���������7���G����u��~����Y��?��#����[���v���R7��gKaT���F�SҼL[o:k���׿���Oh�E�hÕ�i��	��Y�E�&�ɪFT��ƶ�́F�GɽVGf@J�1��
P���X^c���3o�Ԣ,k�	���G�C�����Q��P�g1JF���י߆���m�+�wHlȴ��3�ą����n'�z�ٳ��8�z�<֮���3�J`�F-�v�v�w��)�)���:weF�pQ}1,qkz��mZ0��1s��^��g�|7�)�({�9c`�;}^ 	0�}n���f�	�p/ѫ���C:���.Iϋ�O���z�g�=��.�Pb�g�N,{��Ͽ�xN���,��>^y���`�q���[w�1���L)Y�Y���L=��X^��sRi����jpPWK:�#�c��5V��SU㼅�����x�\Z�4��R�����.��o���=�sN�~~|ɝ��0�צdzA�s����hl�+���}#�F}�kL�p��g�a[�3���wZ�����a�^�����r�|ȓ���$��"'�v�����x�B�ضM�&fWM�,Z��������zj".e���I��H��౦�^g���L%(�Z84$轱���rE�ܐZ��Λק����t	�I�C'ڿ�+w~x*�h"��Eɽ˜qS�zS�HU��cZٝ��G~�ˮ�L��+��g��4Ю�n�F��ǕiMj�������W��K.We�=�R���ܛ[u���{�,O`!@�e��U:p���?�@���$�����:��u���R��Ś-WU.��u��
�&���.A.?ܧ��Q]z�=~LO=����}���o�����$#�P7u`n~���7�nN�ן�;n�����_�:m���ٮ��&�Z���P-�yw�\Hڒe7��M�N�%Hz�z�@׺06�Z�� t�����́bЍ�f�@�ٙ���#��B-5�����caJ[�G�Xb24���NO����V�W*Ƙ=l'�ie�=r)o+E8�njn��k)D9�P�2tk�C,���Yj8m�nHQT���}JBYMkq>�d���}@CyUJU��sY�Ǐu����{��_=���xDt'�<�m�]t�E���n�B���Zg7�Lf.��˿��K�'�o!�7O��(�F�����g�����C��|6�ǷȆ���Aޗީ����
�������E@�畽sU���ϵ�ywU ��o�^���=��i�b�i�G�ç�n�q|"z�>k5��i����4@���3�ˏ�������p|���;1��`��!|?��<�B�d��l�-�{���Gǎεg|��3�4_,Ul]�j�5�9����+>>�9�>0 ۆ8��K.S�\��Q&�6M�T:�_������N�TR=1l�f��������L�8���
Z�H��u3�	:8ev�hd�
�������č��w���k��K.��_���#S�E���1 �Y���`�fI�F�Z8k����X=��B�+�����7��zN��V�_���iMC �T��NґL�yn���/ظ�e�7���D<e���,�H_��S;scI�	��dt����h�_<�cY�yι:x��ecU�m�Qk����y����o���^[]�����xP��[���
��
�T/��Q8R�YP>Z�͛V��3�龻�Лn|��j��Y�Y��&]�XL�;�����J����}1��%	V<�V����H�f���V/�R,(�(��S��T��Q�B�R~K!�i	L�,�* gZ�ߚd�!5�Q5%gRQ-+Fe�j��BiVA$eR��ݝodE�DR�b˜�ꍂ#kE��1��-� �����r��9��Bx�S3�����gs��Ά6L�2��6-R_hV�vYᠪ���f�y���`�Ǔ�|��3f�Ë��h�:�)���*W�Zi�]?������,�����t_�ߏ��Cg!��5OX0|��/ΞeO �?�>�
�ﷳ��p?�]�+��{��t����t��K�±R]�=����9���<h�;m��|7�F� �}�q���Q'��}g�t:s}jLG\o�j}s$kQR�̾'���=�ȶ,���yB������2ubr�.�f�l4�y}^�~	��鉁��S�Z�J���7|l���>l�R6׌�	����_��|�\���hz^��3�<c�����gO�~2�����	?:yb������kh����^^����_�ʹ ���*g����W?��������5��լ�9H��g�āc�qNx����7D������M'UO���wu�@���?~���D?��/�7|����3}��0zә�Xɽ�p�`q��U/+e��a	W�>j$�D��S�e}�ޥ�]�i��>���E=��3����͉	E_v-
6ߊ���Ĥ���:��Q�Q5��?cV��|/]��GFma�����jj�8��-�ͤ�+����krjF�F[�P�\�P��7�b�llR�}Z8��R� ���:Zo��Ơ2TJ�Y8�@+K���yW��Z�+���j�dM0�sj�y�i��V�̔''�ʊ��a��EU�-[��Q!ӌ�{f�מ�����ʳ3���3z��}J�;U��y��m�v,(hUլ��Q��T��R,�g^���D:��\��F'��GT/v!��n6j<������
�F�Bx:;Y\�����ߩhCű�����t�E������:��s�땣
g�P;�R2�Suz�g<�Lf����b�R͢�:G4�蜵˔Nv�y�#J%bnz@a���LU���ėfY�Y� O��}qO�ڼy�\����ϽP��= p�"��F�<(�l��>�L�3�َ��L'�g���W�w?���m���e����7�I���| �����ks�8���<|�o۷o�L�ϰo��������	ք��w��~;O0�!̙�jOn��ZP��>���ؖ���ξ��B�shh��w�Ӈ�:��4Ǐ'z�=�
�Y��͗�پo���ܗ����у�����mO1��g��^K�}���k�+w��*k4��.�~�/�Ï�'�o�.�q��~ �,�V睯���{B)�� hT./���d�=y<*�Y�eI�G�c$�U�[���`&�&���KXB��NEUM���ut�`T���'~�t;t;��ֻ���T����լ�,��q�8w2�_�� ��5���Z��?����w��?�믻Q3?/_�wߏu���[o����Tm[�xp���)]{��&�Hif+ �%@�efjV�.V���zq������ɋڨP"�4z��~E�o�"��
���}KTmq���ߺ��@��
3UsT�p'�5ìw!�:UH_H�2?��yB)F̫E�%"ʥb��T5�V5�*�I��� W7��sr}t{p�J�R��pc�*)���05��}9�&�k�sL��޷��K���ޗu��/�7���z�0��ҳ5C�>�P�VP�U.T���݊�ʊ�ew�zp �xӇ4v��F=-�Z�d�=>�#�#Z�|�ݼ��!X߹��eskkq)��{ �J��j�^Vk�=�Ƚ�Fu��?����zf�a�t���	�Ej�.تJ��B�ؓ��޷a�@IQj��_ǔ�N��i=�{�[}y��f�Bɒ���d'~���|�����'8P���n�j�)� ��݃���������rٴ�&����v=XX�͗ǹ�� &�W�{ )�{b���,l�/�#���BF�6�;�<�d�R�?d�d��4��1�m�-��&0C���!�����>#d������Sn��}t��;���/]��*X�:R�xA;��976@�I2y�������KS9��0��xd����j�%䖓>�������������s��TM8N��["�=���D���+|�[բKG���`ªR�q4�h���K.��o�ԫ&��������I�˔ ��K/����;͔�%�`��>mz�e���W���S#1d�3�(���!!��j2m��bA���!�(� ��N�րb,�X��Ӈ�z�/�~���I�C'�w��������h�_�6���k����i��; ��l�害"��,���������f^Ng�~��>Q�����(���Y�v::r���ƬY�ހ�=�~�{X�Nꐅ��1�a7z8�
�!鼉�ă��ѐ��O+��W8U��p*���2�FT@�-�R��T'<�vV<1;��1"
u�"��n�~w�o�ꡆ�lG�XX�Yԓ�|W��E'%WÓ&bn��D�a	��j16�IZ���&H2Scכ���˨Z�H��JD[J�;j�Nk$Y��>��Z�(���������_�E+7�_٢�߽M;)�V9�Ҹ��k����V��+�[U�̳֪՜���S�]W<�S��ʗ0�̀������#:���T�\%;��g\�=����(�Q� QrJoy�J���ޢ���'�h��>m{n��Zڲ���gԈ�w=�t�Di�h�r���:1傺V�U��u���j7f��?��P�X��dj~̈����z�`���^ޏO<Y�_����3r�B>��G
�Pd;�������,�^ƏG��ٗtMk��-�P���Md8.���ۏq�8n���m�����y9r�m��e�p�D�Y�ξ�W\q������wy���<�}��$㧷�Im��n��6I�NSoz�U�3ӓ��Ojf#Ȗr��՚��~���x͡���x�t��y���K/k�e� �i�!)����6��d42a΍F�ػ��{F� Ol!�{�s�칯����e��|��d[���<�����}�2����ι���J��*쯿�}Ǔ��ꑈ�����x�n��W,;7I�����������J�k�j$�M��ݬ�����3:�(���`.��O�������8��DR�(<�@�g��_�t���I�C'�������߯=Q�t$O�����Q+���p���@�PLAÑ�`%��:G����_�S���V��?���Ol���]ec{�����G�qi�y���Uo|�������֒�sj;�(�GgJ�ţ�g��_�W�Z7��z;P�o�"KT�[��20R���3g��ETi�ͦԠ�˨��R"j�g�xN�hXm��PD�Z� =�����7�hd��	
LN�XĴ̅�8=Y���%��1�8J��г9U�h�����!墮:����^���Q=��ڿw�N;m�.z������?�x�Z���'4�z���ޤ�~�y*LU�R֒���w������?��]�|h�
VV�Z��49v\������ޣv���k�(����K.דϾ����/<M�FB�X��3���k������r�}��o|�Z �����麊���T
�ͧTc=D���ߋ�=.i����J���{�e�]]��7w���=9jFE��l�F�ƀ��=�	Ƙ�M4�2�L4�"!�QB�(�F�������ͷ�nU}o������c�Ƿ>֬�t�����ު�կ�~�}��c�<6��a�`µ<��>��ێ$�BWs�\йxk4̅Z�q�/����"���@��R�t�6��R1�G�_��j��D���'� }�#6I�o�s]��t��$�@�(�T�E[rǽ|0����hkm�֧���`i�ʹu)%U�p����X�jT�|<�Lш�x��ˮ�RP1w�4�4�̩��M���a���LV�iJã6~��(�D�GyX��+˩�a�����]��n�	�_=�{���+�����wD���;�K�ե:.��V�oR��d�u8���O��5VC�P9�Hk�y���^+��5Z��E�:|��[�ow���4G���c��GZv����YG����I���Z��O�^Q%u8�B>��J�|�U8��aܿ�^�ɓ�@�U�F|��b_{IqL�ZvLs�!�$H5��T���uq�`z �e�z���E�.H
��"~�kN9�y��T1��&������G�X2�"q�Ҡ���K���%��E��u
���Xe/�����c�-��y/��Xαy�fxق�'�F���¼���<��s������R�/GP�BrLF,$���֣�
�{�.����L��ֻ�/�<�
M��vn-��P,[�ը!2}�%zY�Ե���m4\�c]����4��Kp@Ғ�9Iw���fwL燠Cw�H]$�+7Ŷ��E26�R1�i�J}=�Ng!��I��,�^�ǧ�}=����A��s.x:�k�����]���`l��~d� �N��{1^�xt�C�sl���L��v�q���������O��ݻ�}�~�>lF_��Wp��Q���ۤ;��<�C8>U��|�c���ʫa��̐���]����v��$�]����������:$�!X���<#��p���^(C	���Ulq��	�Փp�P�ֆ���d�f8��J����[�¨�ԩ*Y
grQ��H���L��w�}��4B�6J��:�Å�N�@���l� h�GC��WQ+l��1e�sLi=�����U�OeC+	J�q!6�l�9�s$�E��s�3�}05��c�g4֌iXҠәQ$᪫���L�?mB_Ejx^
o��C��I�z#� '��E/x!n��GB
�X�N��F,���/��ͷ�c�g�>���)9L��T�uy�����(���ה�Α�'4�ֹ��/�������oI˱�J�FӼ޼.���U*J�%k�Ѕ��x�z|���)��>��خ����!���yL۱L��X�����W�����"����}����ķ�����r��N7Ɵ����̷~�G*y}�RfG�e��7�=����'ٙ�����#lF�8�M����2B�3��/>|�)g?O��*}�RR��O|u��d-�$B���5B�
&���P;�r���礝�ݘ�F��/�����5���-��7����a���{�<�#����
"C�n�]�7Q�5���s�M˅J��d<����733�s.�w�u7"�-��R��O�w�!#T�u
���)��R��E�1042���
�%TM��r߸(��n�ke�d�`p6d爢�4]���W��]��0�"a�����������8pm�ujDsq�@Kf��:Œt��\:Iq����]��l�?������럁����u�����?Ç��+T�1�2��!8��n�����������#e��[aN�(2F�w?,l�͛O��D8q�(j���X�5Y6������DX�n++#)���%�F6�6�]#�E�m���t�ӻ�t��}ᦟ�{?�V����IvqM���I�_�ב��Np�	���+�¹��0u�q8v��};&V�"�&�=.�4\\�tqV����B�J�ϸ 
�:ꊡ�"�w��]�E��r����/A޷
{���Uo[��
�r_�.�"��u�j�4���j%n	1���1�?O�L�jf�X��ف�׿�k���F�Ww�.H���jM������I���+�{�R�:q��y^��Xd�R�H������m���vb��5B�kTk�p���K�}�~�\v)v��-�'Qj�S��� $���������ې��E�B�ӑk��TYN�h�<�G+ ���:X�K�>�=��O#��(��,���pz)QM�*9����7�LK�A)�2�t�T�s����Ě�����\���ԁ�V�9�������6mي��aq��C����^���|w��D�"*�1bk_Ñ��1QF֠Gd�'���c��R8'���r��V/upΰ�_���nk������x�����_�>�8�%�.��
Ru�i�Y�L�9Q�s��,¢�P�\��P8���z�8�k���\��/�wo���/65a��[6c|�:����C�*���=�    IDAT��L��$o6>>��~�BNX�9����1i84�#㫱��G�̋e6P!���E-/��5�	�KLh!�2����������o��>$�.�B��}�}�(o����zH��<	�$&iy�],��Sa���cw�6�q� n��˺�8Q�"
�b�{�$�E���m�`w|dj�x啛p��󇁨�\_�k�K?<���l��	XqA��D6��Yd��Z���}O=s�>��Ʀ��D)�������+�=;Y�,�$�f�-��-�2J����n�� <;A�6�+���]2�};�Nu�l?~r�>���]��9�ބ83��݇$�O��X�fy��*6�qٙ�8kCӇG_����6lX������Z�yf����BaY>Ur��!e`4�j��t.�4ꌒh��7#p�>uõ[jĊ��l
�p{%K�����t� h9�JF6Bn�ƃƐ��85TgE#;n�N�����`_w�!���r;M-�AI���8���{������%GެI[O���ې��P�76�8�G"YD��m�S�+/�V�<':�T~��NN�R����}�Љ4Z-�8�4�}�=��g�N���?�m�OC�ّ� ��:a��v�#�n�P��4~�n�)����/�^G�)گ^�vM�pδ:A�h�_��<o��-hI���^�@J��\��(��mx<�'��q��h���V�B��8��Qc�����ހ� ��"�FR�640(�;99� N�◾w��m{�h�zϠ��F�X�Ol2�Oe ��u��e�w(�!���#0xqOq��'�e~�=e���F2����ə�zT�G�x3
M��Xf%ҠV���u��e 	}x�iZUl�ǆ�<2��췤n;ߗE.�!d$He�fC��*�&Z�����?���֎��2��S'�v�zlߴ'O�]�	��O,�q�9�}�]�=[�
�l�s=Y�,�>�Z��oފ�ax������B��(5ƹ��Dٗ?�*?zXRq�t|��%<�qa�*�C����6\tI�Z+��)�E�Z�Na�EWt����	æ�*9�,�ɢK=h;A~(���DRm I_�ԝw+�,��K�_�+����w �v���0���Ɵ��@�Af�ܾ!��3n�l�ٞD07�U�,,���И9���>S�'�R�XL[5��i>��H�_��������ɱ��+SBHV=�2\��6���W�����h s'��������~�\�(��8#7�$7��������1!wN����f�a��5�~u�/Q��庲����c~qa���Ō��癖��6���ș�������
�rAW)N�h����b��]�h�U���W�T	Z���M�5�+��E�c#�%W4�J���M��
3b�!fnY��8N�D�܉�vy��}��?h��U2o�e)�yXɾ�8h|�R�Ɯ�)�ť�\,:��`����qF����	��N�A>�3q�m?�%O�T�V7m݂c�N`����瞝��K����ˣUo���\����� ����i�?�\)ǁd>^�|>�Ҧϭ:b� �}%]jݽF��L�z�z-O���V'Hu@>������+���������6��f�(ʣ���K�xy���rO�3Y��X�˞u8R�W~yX���Y&�S��r�ҸT��`8o"�hݱ,K4`K{�t�9	�������1ؿm �5��7~�?&g2�QGV`�$�Jw5�<b�I�6x�+Gr���� 8@ǿ���"aΒ��m$m��1�"0B�Q.5�[ux4�	{�8R�M(�ҳ6���Y��"��!_X��ڑa�Or�G�����7��̱��67����5]�嶝~^�'�ŋ��l��:Z�
����9ڍ*�(����ô=<��K�˟݆���G񴫮×�ic'�:%�-zƄ�c�6���"J�֘�S�S=�،�tŠ�9.
�E�T<	m�V��d�D�*&�'���˘�V+��*(6�p�9cx饛p�џ#k�{g,���
��a$�,���`Z}�?�|����?���D�:��F�v�
N���}�ڵn��rm)y"W���Z���b�ք��ю,t"�����5���Sw���GU)#n�/��K7�՗���oE}qZ��� ~p���P�p6#t�`eG�*g#��<�	N	V� �M�uל���^��y8I,5��)�!��HsF&jؤ��g������H�	���4R" ҃��L��r[m��ypn��
�hi���h�4w���_:�T��5�09�e4�1s�WC�c��
��K/��Ⱦz�	���}��S#�eZ���<����c{u����r3�Hul�
y+Hs�鼷e�$�]���I�Ǳa�zqPHj�,�s��\�Zi]�vKS��v�y�R4�j\��r�tI��F�aڦ�F��'��xl~�N����浵���RG&E;��k�@���yֈ[����oe��|�$V�Z��k�F_���4Z1��<�Q�c���q�hy�B��6�ouN�@��"���Z]�I�B�۰_v9v>����<��	1[)��/N�4U"����$ׇk7�a	s�ȿZ�S����	~�O�>�R֧܀~���]}~G3Y�g�ijڛ�κ_�#y�Y��!�ia����4�N`0B',��ȐN8�������"��>�Q 7
��"�|��@Z�:���>�;o�
�,�����q�c�る��v�"�gǙO���} �C���r8x�	i2P�fQ_X(���ذu���w���15u��'�ܫ�+��K���C��āc���^/�g����8����A�y��d��6s�'U���!�cK/�0�)�b�\aЅ�n$��]����p`�i�.�]*��ժ%��z%+��Q���q�[������Ea��=�]|��Y,#��PCe�p�q\����/�z=ra��Q����� ���-7��x/Je����А�ɢ=m:��,!��C����L�����RH��������˰�`W?e~��N<��'�ɖ��N�[~	;ׇ�7op���g}?g�Z�`E����4�q�s�`��=.e�8�w�>d�y!brQ@��V�h���W�Z���FWX��}_45�\��e�޸���¸���oZ�L{n���#��XY���he�+N�r]��o����}�E�HI]�O�,y]'������V؞�Ue2��r�x~+��v%s[s��74#z�7zJK��iB?��1�s���$�9Ȱ���A�ٔ4�\$�8J��yi<��i�"�<��b*�12_�3�8sf�_������M����`2��|Q�D�2�O�k�Y���:篯ܿ�g�~x-�
�G���k�rΝ����:����x���>�_I{i�#����y�4�&
}�pѡra�&9�K�|�?R���:��KE	/��%Âl��ޘ�2=Y�Ԡ�G/z��������B��{�)g?O����o;��~�Ʃw�̠��ty����$�_Ӷ���g8s3��P/8:;d%Gp��h`(c��/��X�Ӎ �3��Y<|�'Q��!�U�i���DrC�ι�M�/
A~�MR�cd\��
�����,U�:mLlZ����@�o�Ҫ���\R<X�52�/�=��E����_q=������#<���a���~�>��Lg��g�I`)�4.MFVt;��g�jF�����"�t��v$��"�#8?#�����XDi�F[��L����\�=��^���A��*�q�Cs�Ovu1�4"�N�6K���e��}o{����$���30;uy?�ُ��o~�b	��cb)$q��Q��e�}8>9�����Ȇ������=9�����mԂTp�����98��OЮV�.��=��� 
�QT�.:�(���~���ܖ��؁Y(�u<��!�ډ�6L�٨b�c�cxlT��T #H�{�'i�h�4��qQb�F�j � �z��'<�p�.�ZE��}*C��U(Z���7�`�4�����O��:�pі�GޣAP�A�n+�K���z�`��L��٨�#�q���$k%?�g����i�xMh��m�Ӗ�܇6fa{V�B���R����r�h��K��/����:�#G���c�3�/5��r>�:�͍0�3T6KK���� ��ν�ed^g��F�)�P�V�y�{Ȏ��{��HW^Q ��Fz%���M:|�s�{S����!5B��h��h���Y1�7�A7V��ޮ5�n�\|ŕ�5��W�8��MB"�O�3]���O3/�Q��RϠ;I$z�a%l����OF�͎�2����L���rb�A���hh�v�J�g��b)	#A��3]?&�D�S���	
f��k���0���x��XJ\L���|l�a�/�
�5�r&�V`t�iȔ�QY��٨a�A8F�ɣ�Pc��E��r���q�Z�ign�{��.���R�`x�*l�t�$#}�����cB&!���<�����g>�s/	>�����,�1|�E�-�Y`8tkR�ݲAg�N��!��m$�#�!�0�R��a���z�r��#`��f���H����3���l�Fvioyߧ�[� ʏ���PZ�[��Rv<�,|�Ul�����#�D�ش��Fg�SG040�k�KY��3�(��1�X�N���80=�_.��� �bM�^��\�+(�S��_߉�rTT��]_����mw!�7���SZ���Ch�����k���]q�D�l�E������i�0�
x�!�:h���J����$�1H	Q
_j�F���ܼ_��rY�F���e��m%�q��[˘��I!`����>���q
���jt�V�»�4V(W���z��fZk�FV#Jux����v
�k�X��J$S����Q"�F�Zʥ�#��(��Ę��t�D�����7+D~���)�2z�/-����6#�	�$-jnW������N�x�;�Q�����ÿW2�Y�@'E�V^Y�zb=4�Zi����ꤤ@5�́�{*�ù��*ܿR�me	����XTd���8<�q-g�6��0؞%�C?Ջ�-�^�W^�<r����	4�ab�t6��A�MGb:a�o�<�6`3�n���2v������9�S�`�����Nֽ�79��R�I�N�M��Ө���-�NӢ�t($�,�oOL�O�D��;A�S���eĪc��v�� qq�������w�S�K�8���	auc�Iʺ�L�kѕR�&�طy����ZQ(�Ȅ�b�UևG��C�������`�i�0�vZ����1�Ç���2�w��h��0���x��`�,".��0�0�	Э�����n��o��$,O��+_S:���C7AX�Ò|Ե�`�����R!��Î:4���>��9
�S�HyS�&>u�m��m�1�(N����0�O�S?����.m>��O�YDҜ����=���ҌtY=v�x�	w;:�nBM�"x0�4Rg�#[B���BY���
VO߾
��1��������~��7��G�#��H�2�Vm�l����QxEOP�Z��VBY��E���K�،���)f`$����!T�d��򘞝�hG�_�ʐh|�E<�d4Z�bͅp9��I�jt�}�_Q!��ѬB�ܿ�y�75)�Xs�܇�4�D�'��\#_������B���Ŗ�P��r[��:
G�����:'�:=�;>�>4��y�ڞ��:F*k�B�$��L�M!�Z]�O5�&
�Lt5���)����R@J��'W��0
G�:IY��Ԙ��
��W2�E:	�AM�V�W�l���2]�|����,H�:'��sI��#��WgDǫ���ҷ��ۨ��`��k���E�k.K�=�
��+Lu��l�&9t��iЍ�i"I �;%�S4+MY0B'��6ͬ%%�*B�4��i�����W�r�)7��fhW���J&��o:1i��{"��E_�t�b� f7#=�-��l�Ii:[�R0����ƻ'�Hر+61d5qZa?������oy;̾a|��7!�q�y�������|	�sX�v>~A;�K����� �N�VN��}�o ��/���2WM�ىP]ja��3q���х*"/ۣ~1q�t���g\�m�7"��8x���=0�G&��<ะ�r7�%,n ��B:��X���db�&�=�z�8t�M($	���4oڬ��Ho��M���4ј9��?�<�㛟����[1s�Qt[54[\�������w"Dd��et*�x��O=�����}D�?-lY;�N0W��l/�t���DL̲s�De�8z|��2���[�z�F�����#��K�{��W������_�����W?������I [@y|f������֕mt�K��͔p|��z����V/��č�0�:"����<��b������0͔���0F�8v�k-��5�-Jl�h���/�(�"��R%=�"��s�Z�?_��x���ꔧ�i��1p�g�@�J�,�D����B�JD����5@J��o5
���2�v{����҈k�^�o~�y{�_Iw��%�퉴�?��Q-N��ЍD�p�gj������c�����W*/�5�U�F���h��f�7m����\٠�q���s��U��S�,w��5/�f�4M��3u�:�cH-���%��{��]�#
ݞs�����WGL�q��'���Դ ǿ<.��1b*�I�j^�Wk8㬳��<?�u_����0bv�d?(_:V�4�2�fJ��A'{��8F�4��I�n�ǆb�{��5���<���2ؿ�8wԓ�7��7f��X��b�):@�μ%Vt�Q�����f��#��P�7մ� ��R� f��YJha<��fe�����������b9�����w��y�a^���P7�C�9��GuZR.�2pz�$�yso&�m\������)��6P�@�)��3hR��y�(�1L�(UO%=��H�>�u�@�(�k��d�L��;�<H�$�I�d��4hSU�pwMt�S�;��t���o�L��CDT�#|k��\{��*x��A��?����W�0?yc�Cx�5�Ɨ~���K0G&��Z(g�1t/�������.�j���0i���������G��_16�V#����ѱaY\����/|N������e�������7�O�zl?�������,��,F7`��!��e�����GhN���X��;��5�=�)8xl���/�7��KKضy��Q9y�mǚmgc�����0�!t�x��EѮ��4����8x� ��D~����t�S]t��U���ф+���H`�nT��^4K#����s9Y�5W�Z�9�W�W}��<�������Z��J,S❔�!�g���Ө(�]����<��r_�^	lZ���o��L�+�'E.4-�\���_:!�l���F&���c��ݴ��Q:σ|�2ş�<'���q��\2�G2)��q(iM)�Wϋ���W�� &s���4_M�ι�<��US!Jr�X"���k�++Jϑ�t
��p9�+��<S�֭�n�?<'��z�����uP&�GQ΍���p��G�D��N�F.SD�q1;=�g��k��:�r�1|����gV�R%��iйpz�+�c#qh(�m&�H�c�
��!w�лv )��������܀~���]}~O#���8=i��A�{#�	537���G�ʉ�c�
ѪW�-8�<,3����:�9�0�&���C8q �h�Tp�P����-$$9d�sG�̻!F�3Q.e�\�{�o��;Di ן�MРS�Z�:�aXn��j�I����FG����=E��e�aRDI�=�$[@bS�j,a�S]
�,)g��L"eki�F��&s44�e��%0]B�0wL�AV$O#;�L���md<Cڙ��y���g�O��j��y�L�.#;�w���_h!,�~�,$���^����y�w�lXU��5C� �1c��Ww���z��ߍ�ŘL�l��Em|�_a�o��l?[w��g]}���_��� j� �⨔�e�U��C�z^s�8~�����7�t����� ٛ    IDAT���#S5�4C`��q���W��g>o��w�k��	��u����7& ��v�I$�*r���܇����� F�����5[i֑F�+����2�����Q��Q5�_��B�گ��s�Ş��_:\Ե��>�U�3��KIsRE���~�Pi�W#~%O)\�s�]�5��I���Y��/:�*�Ks��ki��A�����?�E�Ĩ'������'}�{�;Y%��Њ���L��hN�J�z�֚�T'E`�[!s:�C6Ov�/��"u(Xſ9�:GJ(K#�4���5�D*�2B���89�XI��A�}�y���'Z���X��.ǣMu&5w�����zp�`(����&F�H��\;�1�T���^z�+pp)��z:�
�"b�GfWZ�R�Z��^&(�C��B��
�/�&�D;a)p�#^��\�d?�ߕA��z��k��k��s4�5#+�(q�ä0+xQD���HB؍
6��<�H�C&�k��6Š�YIf7��a~ҖZaj�G�/��MCld`D�� 3j#`��gG��D�ło؈�/#��f�!�D(Qt��ұ�JB��x}����@�*B1XԈ���!�l�ȧ�"�al�e�07n1wF��}��W�fK��E� �a���`:!����R��	/�<����%���c�Ab�pa�-��)��i�B"9�N+A��d���b0lwg�ss��0�F��w1ul����G}iFz�S�n��a��tV��(��I˂�t���5��|-���z�p0<:����4�LHs�v���B���G�-���GE?�����T��-��`l�cv7��p�UW��a��k,�)"�����TN��k�7����b|ըth#)097�T.t�;�u�*��)11��U,��Ԅ��S�����= "4=2�W^�i���k��m��$+��9���eĨeW�W��q�d;+�ۨAѨLIZ�j���05�� (T��;�?�SN��Q���4��WgI�i����!��e`⼘i���]I_̅�<�8+M��^$���d=O>����o���{HSiI:kz`Q	c�j�+�������}Q��d�:gz�E��Ө���Ы��7�^wq���e��)"���<	���r(�O���:�~P���)\��	�Z���X�.��\v��f�7n���!�6-���$B�j�a�K�,E���+�OILf{$:�F�R�n&���fl��_�ix
�����Ÿ����C�>?�J�e:��"�h�	<�V9k#�Z�h_AF�A�F�.@8VA�e��'�42]��m��mɻ!����!3�5�i?eZ;��O�0@T�	���2D�Li�J#C����7;Id�|F�9��X��̞�A���mG',nS�3�a��.+	m4�4�"C�ÎӞ��KW�p�|�s��\�t�t��+:�3���?n���;�b� d���A�\FX���0i�cd���iyX�Y0�^v.Po̡ծK����S_B�711���чatB`�ad%Kz�7�s+�:,J��))���]������fN_?\p%+���<�d������ȑNy�n>{��G%I1���mϣ�_B��E�E'���i��tq����8g�F�NOb��(��$͓�f�h5�ˋ4jUÙ.�i$�Q����Prq�5䂭�F皧ըM�L����.|7�7揪���T��2����4�l��$�s�4~�F�H���2�Sa��V8��pE����eĻ� ��]#��\{+e`+�O��J���yl��9���#ZD�V��+ɪTdIZ� J��!�B����:�����H���~�䳕�B�<���Q�|��q{��:�B�����q����Ou
�I�{
�+�g^��p[%��s��5?�����3�q��|�J�Sނ:2�\Q]�]�r[���)@
��}�q�&\�c�b7|��s�a�.|:4�t�cgC>�D���A�J\^')1N`y\K���c��k_��t#%�"�'�o��ZJʯ��O��b�?�
���@ca�G���;v#���vO.��ci����c�K��BJ�� �A�I"��C?IR�a�΄�CCb�Y��r�M�zy���dK9t������%2�[;p��X�L.���fNJۜ؄Չ��GyV;�E-qVcA��\<��i��S3��l�b\L���;�{<!�Fd�"�9�H�⃑��H�� d`���1,F�1�(��#�!��:�ܒ'A^D!�IN6#�BH�b��D-I��m�ZM����I��(&�a�+��#��zK��=�ݐ%.y9�(�^a���G�h�0�o3,���X���v(6c���D3`^$B�0 �S�[HD��J2�F�c lHz$�m�N	a%@1i�9��nOb���l����0mW�+�L�p{��Ј�"K�G�W����¦���홓��mJi�ՠА(󛑘��ѭ��U�K��Q��iD5��W!m��jĕ9-F�JǮџ���ѕ}��X#5�Щ���H�Y$Q�7.�J�Z�H���C>����y���n���K�-���1G��E�):�~;���3*ƃ%}^J6�A��G�4�QgF/�V�D��9p��Y������<w����)�OS�c���\7e����[����R�J?S��ekZ5���U�H��n���F[��S-�֠sC'���v<���
�����dؖ�)�ܫ5lݶW^}�̅��oލ����EȒB7A����GJ�$�/G�R1�'�k�
����o�����9E^O��p!~���7|�>i�����+��\-��g�8@эQF k�(���a�y����Z�w��aK��{���=�QL�\�(�6E�X�ż4u�-�m
���E�Ƴ	�D�6��,�Q�LC� �rm�}�,Vf�����[w���P���.���!0�g�&���	Y��QQlA���v�~��e�4/�H���4�N]d��� O:U�$��P���?�X��:$�[t\BX��Mb�1��#�,�\�҆%�bJ��N�bv1��Y��r�,�������q�,�1��I��:2IK����.or�a��������	빈�,fl�C��μ\#�ɣ���02'+U^�ʇ6"t�?4����Dw~�&eMݸ-�!K�r�2�^���,��@�E�����(���+���ѩ�,G�-s�M	U����%�=�}s᧎���)aLET.UC�q͟,�w�e>5߹Ұh����+�k��)���z�C#U7�"S�Vsۚ���Ks�J��HSs%[\���������h��4@
Yk���C�:����0(J �'(�����4�M!d۶��k:CIyA�à�k�5?�i�>B@M�e��ֲ���?4���/-��,1�'4����>�\;%m��ثQ��@;ͯ˵�E��s޸�:[�8p;�C�;�:S�p|�ǿi�v
�w;)��m���+S�Nہs�z&�>���d'-%��~RL���8>$�e�+%�1b�A���d�h+'���>����}O4Ҝ�)�zҠ��q�\R|�G�X�R\�wb�,E�M�Ag^����������mB�T�I?ħn�sm�y�-�FT����0ޜ�$�<��2��96��jl�)�,���i�ts�
��h��\�fcq��-#�q� ������4���z>���ý�����@��e*��>K7���f,�v�J`�vݰ�;y��YO�aw��x��W�!O�<���t�b�4g����M�9trH��a��nQ��4�L:�5o𸀗)�.�����A����4&��e�p:		��@��2�g&	b�!�S�2p�B�ŖsJB���|�-:S�Q���M#M�%�`�C]l'��� �m"�пq�	��.ΞamQ0'bs�q�:SiϗV�Lo�k,�*�~zngC�v�zK������-tua�A��Ѕ;e'��#���(́3��@�Uj^�zU��U�U�+1���:l-��f�ra�MF�Hp��x��iKR��r��hU!W5�+�jD�R��C���羵-��w{e_yJ����,�7���|j�+E4�!9�^�A>�y��9�AD�G
l�I��-G�J;��:㩓���"��Wj@S��}+""�n#u����h�a�q쵠]ITȝ��Dkx|-��{H��2�/9Kr{%��$����7�/�[��
��z��0�J��h�]��+���K�K���ȆQ��`�E��^��Wc�.�_n~kX�D>�JĠ�g���J���ז��2D��13y�C'��!s�����?`�9�S���A��9��������1�q�y�t�7$����v"�-��B��};�����f��-��(��O�
|D��ЁC��x��6�T�Ƽ�xS�p��f ��=S�u�NTG�� j
/��B��^}>n�ćq��<�� ����'̲t�
��~%�d*:2ا]4��Y��CML��j�a��8Y�Μx�M�g�N��H�`ގ��0}@�IX�mV�e�N(ڰi�)�B���B����29T�!lfC�n��<��7�����\x��Xhw�;Y������Ё�4�	�Q���D�!Y�!�x�ST E,�G���߳�bBۼ��*`����k"�,���6�9~<�`Ď�3YW`��_&�i�]���ad=Y,��O��>����L�3>�Šo�[��rF��G~ ]�Hr�����$2),�D*
��~R�T�F��Q��m5�����8���,b���5R4 -%R���E��ʡywB���<8�#�D!o��y|��5��\�|����U�F��>�:^=Gݗ�O'YE��64�+#t�K#eqJۊ~J.�s'.�]x�����8:G�y�iX%�|�k׭�2J�����H���p�F��>�Fsݼ6$��=:J������uk6�r7-E�:��ܗv��oq6�e���a���rE�׼���R�qW�D!w^����HMAh���D��3�%]d���������o����_kt���U1 Ny��!��zڃB�f��pr�A��b8ii�F�4��7�M|��׏>}̘=El��I�����F2v�[��d�o=jI�Ox��Zi�p0�*���`G!�3֯F�Y�C�c��`�O`$��Q�$����]Pm��M؀��d�#����+#�ŴC��</+pp��CGhth�XqUZ�^}�K�o�~;�V}��	���xޫ�����w�D3��Z��w�1w@��|����]�,c��*� ��,!\��ad�<3B�pe���MhĠ'��nkf�J�/��5��������� �m�؜z�!��
�%7�Y���:�6��0\���'��lἧ]�G��ڳ/§�}�,��J��C����$lP� �WExBچ��DGD\sZ�8M5��J�`	g!H�/�*%��A�d�tFn�exp�y\�=���!�]C���~��Oc�c!7z>M�8L�hP�smVc����V��*�s�X��r� �88�05s�B@�0Mj��¹�ŊH�Ֆ%�/���O�K�B��/���Fj*�"�� I�B,yWr����ZP�9�c��x�e�ҷ4Ϻk6!Q�Μ�J���D������,h�Z�k�3���8�ǚ��P�� �|�D�9iKU%�cz%J��P��N�o�Gamurx栵����e[�� 5 
�9���/��:���H���|r;����RY�|��իQ��{��t,��؆8U��e��>��	A d��B�<ثdH���Q/�'G��}�����)qԕ�p�6��6iڌk�B��V�j6�z:gt�Y�ɠ��'ޗi5@��i7�S���4�6�/�7
��v�4G�j��r��4��{1E� ��+�x�u,q��lSӓ��H�sۃa��z��X{���}shXC�7N�KɃ��S�����<y��Ƶ"y^;���\���7�r͕��O�SiV�����v�m�v�U3-�_��?\:v?�>ՅȨN�+#�Ar.	Y#�������'�S�V`��z��3�u!��1�am��۵��N�4��6�v�R�ss�P�r���+�5BDA�!�*�p��ӓ�6��7��B��b�W"ʏ`��7�H��=t��(И'�(u0�����}h����D�su�cW�a�ɼ0���)��T�F�0��H:r����k�ek4�����a�z�N�(/�/(χ�UmÇՐMj��3p����U��{��X�������b�y����^�'o�7�����=&٥��#�D'��e.�A���f��F��K�ώ�Bzd���3�M�BĘS�=c�o4a��g��K�K��y+.;w#~����о�ؿ� 6m?߼�x��7}�A[��d��
Et�u��^���]�]��2��;��i��XBmn/�W�$�}�~g����<�*�s9�_��\sV�Y��}�BQ�;�?����clha��nHE�lIX$1��׏+��Bt��>��=���e�p��f"�����KA�O�믿^D�G�vB����}BȊ4�b������<t>����/�bH�\z1z�!����G.���h�U.��jaӆ8>9������s3�_����w�X�j_��Wqr��M	��8b�ڝFW����i��^�r?�&��-�qo޲���w173/ʉ�N�,-�d.7�������x׻ߋm۶��L�=F�������ǎ[n[��&�5k��?���?�QeޚR��3S�����-o~ffz�X��G���˻ص�Q|�C�$�KK���{���_�T���oÑÇ��R��cR��_��g?���P�c��P���^���U�}5&������'O�m�R�s�����|��ԧ�j����f��D��+������T�!ǂ����۴��8��?����k8|t��,\�kd�w��-x���ajrF������h�����m�{��.~�� �ͣ�D��&Oƫ^�J�욗����HȻ�ׇ7���p��^���Ƞ��Q���_�{�2�j9�=o92�N�:t��T,�#�.��p!�����X'[@���8w��߽�V_<dL�J����=I��{��~�С��n��hz�����8�:�n�u�NgU��Z�w��z�^hu|sa���[��Ӟ�W��[pl)ď���-����?[���`��E&}H��a�6tuI���D�n�gg$J�2�g-��t�p��z%-q,a�KI\����M����n��8+mYq�+g�V*�P�.I�g�1��,2=��ɼ[b#�7��M8<WGf`ͮ���Ŭ� ��*6����s�b����΍_������d�ƣSK���KH:1S��"ܜ�C%�N���u��D�Rȝ� _�G9E����D����zC��sة�N�QXD�1��l���e�������[o�Y����m[�o݌����������ڏ��G�����J�/6}OƕaB֔InO`b2��	H��zA{Q��LDݔ̔Hu��}�	s�@ �~7}��m�q�������֭[Q�����x��x>���c�� r�H�c�͖D�֨#�)���0B�KX7��c�`nr/r��R&����o�(��b>'�2>6��}�s������:S[7n��[�
��{��P���Re->�����|��o�#�v-�<׭]�K.�SS'� ��.�i���[g�q>������������{�����/���Ӻe��#�W}�Y��ӟ�7|���N�o��oߎ��~6����c��@��J��i��:㌳p�wo��is 3A�>���?^pI�;�@��G>SJ��qC�l�����6�}�8~��shx�B	�]v��)��&�P�1�,.��<��U�x�;�&-��	�"n㵯}���r;vD:�)C��+#O��+u|�đ#G�șbFv����Mر�L���s��gS��W����x���G����I�$��hW��=������Ȯ��+��u�M��*w�/�����;�jWS�?���m|鋟���w/���O۫��Oٶm������\�R)�H799�k�M��    IDAT�����{a����	U��.�%���'f���	t�D�l�n�Z|�S���G�����c�Z���
R�?11��S���}LВ\����
�ܱo}�[P_j������(���{vc��w!h�0=�B��#�_�iO{�c#U"X�-�]����$|�%H��p"3��&�֦a7D!���v��qѸ���˗��]|r��ա���?�o߾��ٳǢF0a̓	�'I�.=Q7�ME1H+Bެ_�	/~�+p|����1@ma�aɐ��o!a���rO����>֐6�5x�#2���ͅ��K��r�)I�kz����A6�A�K�-R��,������C��?�����
b�ٿ�ݬ�C!�Ln� @yx�����v>���A�o�k����N��mǅgl�p�����}��A\��Wb�\{gk����c.��ш9B%��j�\~�Ҡ�Ab��i��[�;1�tjȚ�n���Z�g,�������v����"4��N?"/F�g_p������`x�Xn���-�*Yᵦ�=u�}����(�YbA�U(��wa��T����%��ȸ<�;�!i����Ř�t
*��o�sd�{}L�ջ(z�~�u�w���Az��L�M���r�@;H�
"�-;��<�oH�N߶
a�(N�؃�OF���]�l��lK��O��*����`��Q(`��-8x�܇�׮���eΆG�Pi�%|�j�C4���D�JL�����O��)��Ib���AP�����a���Eb�Q.a�j��k���\N���$�1
KS39��#��λ�^��	|��k~O��o�^���$���w�Z���>�l#Z��9�7���2�~x��ၒD��O��6"/��|�,���<���3\x�x��!~W�L��2��H��
Q���/�$SoB��[x������\��M�� �j�LN��ĉ��a}V�\x�y��_�B"/M$�7��Ȫ����w��	�jb�ڒ��^���ྜྷ��]��&J�`��T.wp`5���//F�ͦ�|���.>��s��ڛ2�U��0�18W����Sm���q�{�9�>yR���ڄ6Z�8C#Ø:A����e\��H:^p��ػ�1A˘]��H�uKh�}8.Q�&:$铌�gp�q�w�S0=5+�Q1�C��/����w=�S�L�1�W����,�47�DˆS��}΢V�8�'bT�~�����!�ٷ�d�+S�N��6!����Ň����3F�\<E^�WE��|��}��2��s�N�b1н����;c���[��/D�n"�;!�ȿ��ο#c�����=�`phX���r�u� hV�ܢ���f�&㗆�P%!�������0HTa��(��T��)�:��|B��v�R@ǲX�%,.,,��$C��o�ND>�ɠD�	kR��]ʘ;$�X�R�)#q'��nY�6��~֬��Q�� �A׼�8��>ԗ��2���أ"�09@�=Щ��N&5�q����/Co��2~G�𻦴��]zڹ�d<�o#l�b(�ۋ��Y����<�r�s�ibH�f�CŚ}
��Ѩ�Q���hEXj�X\j�����o�C6����az���� �K��	2}�);=h ��IN�͒����eQ[�K.8�E���ȇ�F9n�|�@�
��,�g'�����0��̧#_�f|}/��#+�iLNV��]�/�ar�,V�q^�Y=���nY�&⨃������:�����H<G򹅡1�l5KD�N�`�Bq N@��p�lŉS�×��G'4_̡M���Rz�o�?2O�z͚^�vk׮(�Y�V멺��o��ƞ۬eQ(�i�F���|PZ���8q|�,�aV����v���2s��KP�5p��Q��������s9a'�p�ۮ�c�_2��ž"֮وf��f����~�<�(�&A�l+���A�N�������r��������U/S=�=��al�1��Z^��'��R�G���BM(!�PBӋ)�+�ظ�=㩒F]��J���O"~�{���zY�o��"�g4*���9��RQE�&��8UP >7�����0O��s��@�b�Ĭ%��P �G�D&���rss#�-[!;f��|�Y]�vwd$1���FsSƏ�u�����_�lJ%�v��s��?
�Y�˰9�x|�3a�8|��h��:��؅"��(�s�y� �7���N6�&g����1�_}�Z�t�K�6�{*�*?%��e˚��3�"�@6�^l�܅X8"ʐ�MD7 i�DXx�z�aUT��cLg���=���<�ҵ�xBj�ۄ���Q�J��9�\AKSƌ��p2KhD#~ɞ߲�G�������+H��삍�W��I;�4��t��	��u���A�X�W��䵥����T���rƈC�ǋt���<活q�ŧ�����Mj�����̿�\z��Յ��I9��޷��:D'�MY(�h"!�2�pk.�NIҫv�e7��^x����,�$��M��'�AՐBɋ�yD+R�$&N��M�6I�OBM]�i�9r���,���ї�*1XE�=������HCӕ�DCC�� <D9�mشY<�0��֖�`ug)6|v�Jv�}7���b+5�d��!�p�ܬj���;�mM1|�z=2��9+{-�l-_�m��r�;��2��ܙr�N�;	3꒪ꪠ���΁����]c1��g[��p[(o��	m�r޹�k�2��p�Ne�y#rf�tg�P(����߭�Fke�pg��O?�E������` U@�q���ry�2�z�*}܄q�8���Y0)����5��E�(�WN#�*���!�a��Ł�q����h�ƎP+,�CX��zR,�voºuk���Uؼ�%ǅ`�%�F"UD~T��;�^-�/�.�^*adc�~~֭_���"��L�.|�����K.���A ���H��$�1<��.3g��C��kVɮ�)�BҚ0a���xe�[hi���uժU3f�4��7tc��do<44�ԍ���q�)���ۘ4a�pG��q�礗�'� M�:Y��$Oދ�z[�G����'�aĈa!�Y�Zv�l"g��L�4E�Ƭ�lTyO�^��݃e+��������`ƌ�X���qy�^�֎�k6�jC��B�M#��W������� �0y)cG����hݴi�0z��o%uD�-9r,� ]]]�ho�霄U�x|m�8�10�/HDb8)\�H�3f�^~	[�t��y��t���_wO�L��s,���������$"Q?�L��������1�]`~��Hw[��1vl;;�@i�qE�#0@����Ͼ���w��o������#:���m�Y�i�l�����p���/�ߛ?\�hc���B�� �xsfO�^{����#�����;a��~���ۘ4i�j���P6�B.��QG.뉁�^i�|�(�qr��X�l1^��v�q*ҩ��!S����'?�	:Ǵ�����A-���x��X��kL�1��)�p�lJ��ʐ�V.v�?au�{yx���� �?$ʩ�+��t�9̩/0��a��_�Ҿk���_�[���S���t�զ���W��'��M�@XP��:;�T���ԌB>��
��>:�ND�\�ց!�;��T�=���{A]�s5�7^��M�"�>��n�֭J�K��k>'��#@�a��Ue�+O�ҏZ����W��|,t��Je)&��Uذ����Ր	�L�&O��w�zCr�$Q���t� O�N� Z�"�LT�f�}8�\��YhT���_��,�(:�	��[��*BU�=Y�$��Gf8w���f�c���'�$��(ጟ��+�-��z6o��ٲ*�lxL/�n2jрƖfij$�q��U�k"!ͱ��/>���$�E��H[p� �./�@Z�ph�G5�ZQ�W��º�\�����a��q[����oF����O>��NA�`K1�L����~����������Jn���8�n�����>[��+�ƚ��a���>/®��(����������n4}8����k�Q��^��qEp#�h�/P`8����vp`@&�D� �O������+�K�G��56�, ｿ@����D��E��y��+W��+���X$_{�59E��Q�(	�|ܝf�1c� =���f��K��u�\3.���!�{�;�Nn;N�.�2"4�z��s礷ac6tmR�����:j�U��]�blg�|ӥ�PQF*����bي����A8S%����D��TO�8?w�
����䆯{�������g��s��b�_l��`C�)�'��ɽ��9V�����ދL�&K��F`��;���=�p(&��ԥ����B%��wT�>,�Kć�9v4��s��8�^��f�9�4=r^yu��͘|�� �"�ZoΜ9Ҽ|���9p���a�ԩ��e�8�ee|��0���M�c�¤	���/�c��*�k`�ٳ���ﾷ nC��Ґ���"���q��Ǌb�O��e�D*��QG��+�bɒ%hllA&��?�[��6>� �5�t
�hChj�q�,Z���l�+@p�t�~��x앏Q�M�<A���J�n��� �^�V4�*E�~C\<5���f9��ZM�����ڰ=��Xߩ���G�-Y�,�dJ�6�(,ܼq'��ʲ;�M�&�Ԟ�]���vA���l퇇����\̉['9��JS���A�U�(�-D}}GC2�Q^Q7�-&��+U�<�c��%1J1�*�8��І��tf"<@��ed.�	Y鰜2�MHg�ԍ� d�fIԣWjѨ��iP�4dJyt�j�Gw�ds�Q�ǂѓ��e�`�5�܌�4��H�+�q��Miۂ��>�4�#���Z()��v��P��"�RZbb�����
�p����l�ɆS9�7^_P�c��%;���
J�ܷҚ
��i#R5���	��Ĳ��W]�e_�B�N$2�B����0~�(�sذ�+94f�6Y�&��G�8�5�Њ���v�q\r��8p����Ɏ����Oi�P��u	3Nq�U�����sત�w+�6�ॗ^¢ŋ��>��&l��Cɮbƌ��>m,֬Z�xO�>�D�(	L�X�˴~͊�e$� *�
6��4�bW�� ���LE����p<_0 �V0�&��2�G���[�6����Mj�a3ł��c�-٪����녹�D�$+�(t�ˡ��#�y��V�m�a�ņ���H�رc��U���Q�ڈG�)Lm6��_�3ǉ���#Zư�Unh�9[��[�+שU�DJ�3�4lV�<�9���R;G
��0Cv�@��R8%���*��c��I :5�bmZ����L�� ��V������ɹ��$�kb|S.��E+�@P�Bх��1�7d}�J�5��g���M�?�U嚢o��*WY>Z�L٬�8IS&I�X$"Ϗ?#Ɉ7Uvx�˵Ϝ�{ѶL����k�5S�I⊂DU�ŇSC�����-M8�=0}��.?e�5�{��U�^�s�Uz|��^�<U'�?v*::' ǚjǨYG�����3Bc���XQs$�E,r����"c�@V����S�S��}�;%������8j�Ԉk�Z�����
�_�˖���N� y���W����'�$/jNC�R$�y��r�����K���#G��/b��8��3�#��^�,��Yx@)�Mf�+{���w��T��VWB<*F\l�Q럚�	wrJ#L��L�	I:�7�GG5��<�}�BQN���}�_[��\�E�;�:�/0�`@�!^/������_(�Y�����F߰����o8׉�V�U���s��q�Nv([A'i�@��Ъ�jI�ParZq!;����=�wWѹoټAn~2�I�aAc�#���Z�&��5a�g�	��	�R;,xP*�Ne�1a�8�>�Y�W]��x���ҁ"�l\F�'O��K?@�� ^v��+����d��|(�Cn`#N9�\r�E;a*���$4�LgInr�幋C�F8�h:���q���.R"7+��U0?}ҩ$^{�e<��_`�M��M�l�JE��� ����U-
��R����/�` "�
5�T�%�*f&n�	�ͨ�Z"���U��e==�����W�)m5�O��������68�?��\(�ȫ�h�C�I! R$�gn���.P2�t�"�%����(��$�������ך��
y+|�;;��b��`aL�⫂�C�D-9�pޛn8L�3uYl��-͢�,h�V�p*L�v*;��b�(�{�"�BbD�[�/�| z�{���Q�4��OkJ�ɴbPF����A'�HE�����4��T�ʤ� �e1.�G�l��.q\-l޲�&[��\�5lnY�y����I��J�蠘�C�:s>���|�yE��1��Υ3���̆��kF(*�������M?6�Ld���k�D�UT��-74���Uy}~_D
�pjP%W橷w�5Ân���4u�Z,��ѡ�W=\t��J.�U:e[H��H�/j��xe�f�2<>L���૯��H���W������R't�ca�&7���=�4�>ٞ�_}��TA��G7f����{N��:9M�����U ڲ�s�$(���hY���C����"�FW��LX���m�4�$�1T����,U�R�ሇ`]��ώ�+}�����2+�	�6q��8��F&,V�x5�.�L�x���U�8�f��C����	�h�g�}J�-Xdm+C���oz�S�]ݽ8�����/1\�QrH1U<M�
��OD����$�EIKRQ�k���� d�@17 '?�� �Ξ"2��k7���+w*�@8$0�@<!!�2��,ښ"퀲7�G����H(/��}D��[6����b��5ho���,�UƎ���,[�;L��c:����(:B����ѷ�s������.C��	��i!�5^HgU������"��T� -T4xL�����~Ր\���D�������[~�l��l��G��.��M�h����l~�Y��v��m$��ѵy-�!z����0}(i���B�~6�����5@�N�����H�u˘ղ%�k��f���w``@�[,\�E�f���u�Q�V�y��P8 ���P�SdcMM
�Y�����و�i��%�G4�C\k�_|���GX��Bn=���(�Z �a揇�r/@sk�ɗ��?.;]��JV�&OB"�B*K��4ze� Mq��k=�F(�s!�R�ƚ�^̓�ϕ��$X����qӤ�@1W��ה���(}ӆ������ ��Gc y��>����#� ]LB񔋪��g�(eX�=�ݑ�6|nl�SC�t���P4"���y�[�-�v��>��f�E4�<u5hxJ�.VQ�F��u�ɚ!U.��	sS��3� ���D�tz��Oy�S �CE������VhjG2�B.��7@ �p.���b���X�t��dxͺ<(!��]���h�� �.�7*�lG�n�>��w쎨Yܴ��/��ǲ[L�u�x�n#]w��Ex{��w��?���D2��믿.��zN���T;�g
>R�Q8��M�8C��t`ƌx��6�Ɲ����@��J��m.���%? B�2E�jb�[7�o2eY3^�M&u���j�:N��]��VKl����u�tqW"�T�M�q���!�1z4f�bp��]Qݿ��}��Q��`�	"Q�J��#��W�[�TQ��P�츙��0ޠ)M���Λ��0!0��u�)��'a�c��u���K؄�~u.8�"�۸f=��h��P,��}nj�bk�V,]�3f�BS#	:�y�S1O�r%/�>��r�"�D&d�851O�0N��� g��,��:�D2�a�"�|��A�_2����J�ީ'��n�	�pH�F��=/��|#��0t�L<�9]��ɗx��S��$*
K!	��Ȧ���� �SO=�n�C���v$�t�,9~q���-��\f��C�,ɣ��*�3�E8����l��M�b�%�1>O�? ��,Xt��    IDAT.cX���_�u{�zp���UV��H�\U��%�/iz��:��&��#�����4G5d�ׯ4�t[���}�d�p{��H��I�QE�G��U1Qu��\	��<<Z
%GH�lHvb,	k���ɤ;�o��X�L	E˄��)�Mj�R�=�Is%��b��,m�Se$�B=�_��Yxt�3:(
�՘hX����'��/��e-AP5EDY4I�5���zE<+����w��)�_E^%����������u�!�p���jA���'B��5?�QX*���)�r�Ӥ�ou�f�� D��5W���Qgdٖs���]� "�L_�S"�6DN�jM�'X%*4��j�i��)x�rȉ܃��V�)3dcOΛ��7���1:���)9T3I����0a�75��X�II��Ux��Xw#������\w�	�{�Ǎ�D��ݿ��w��?��'��3�z�-a���v*��/C��Ö]�x	.���H�a�.��m�2����H���Ԥ"y��|f��K����7�R�P(v��bѨ�=s��XJ��e��"�nR�~���;����;(J~怓|$�k�n�&\��P_̓���5�6��.���`7��֊�I�8D��`�}ƂE_ �#�Jr�%� OR�V�k� �^]7�>]R�Xx+0h�I���P>��"�:��}q�ݷJ�I*�4����~{կq����w����%�I�	8�ԹX�ѧX�d�q��iq�*�5MwE�Tr�
��&���-�����k�1f�e		��#��,��]@ȯ��<�׍	cF��'�ES��+Ul����c���Fv8���(�#Q%e*��%�'���I��҈�M�)D*r���L��U@8�!
���[o�=���mcTN��Y'�� s�,;���8Lf��,��b"� ~�8����5X��-�1͐}#��C������y��D��k�ŞdK3fp���b?�k������r�d��	�>I֯m6��k[,D��?^�m$�2IJ(��76�wr2��]"5"�!]a�G?�f>XYG4��`cF5b���(fm�0i��Ia�{|n���T<'M�۬"���ߠ��B��$G2�\�[W�q�U���K_̆*r��@�wy�X��/���W�А'�v�\�:-���	#��$��aA�
Œ�nS�����*�3�{B�
�>ғBbl�yE���y���Z�Y,Pۈڸ݂��h��F8���)>��y�j����lu]B��>����H�*�"JE��Hd%zF0��?i�Dq*�5�Q�W��R%���JH$��s�*h�gx10jq���*��>�ֆ�E�j����<��p�8��X��x ��1gBGխ�T��'�D�
�G�ZL���v!�M"Qua-|�ZELo����Nʷ:���G�K�j��O�]���x/���'���s�x�l�J���� ����-�,%.L2�b�,9�ӈ�s�8ш>�ȣ�*B��"�����$����:2�^���YgK���R����Q��"�w�2�+dA٨�&�5Ne�m���gr�\���L��K&4���[egI=:Â�H�~�4� ̥��y��pR��w�.���0�$K[��9%T�>$�x�a1h�͟��<2�i�pv�g ���!�3�1�L����=�g�Y�f�&��֐DLn��f�w�9x��1u��=�|��]<�����+�W^~�_��}<{� ZGvȁ���k���-<Ʌ
d�8�}���y��b9��ވL�F2��O"!5�~W��A9��3O>��g�=B��9Xa�n݌-�c߽� ��}|@X����}QqU��/`���E{�h9$	s��d�M&��U��i��8i4Ƃj��1����p�
�#m�:>8�VT��*e�p=�7z��Egy4���E1��U��V��O3����q��	�i�W��R��&�06����V�$��z���6��-�}&Z�:�&џ���?�h�k�_��ŇwTK�Z�+(�E��H�Ěu2�^$e��T�,�����D@M#��\��f�gx�J���q�A���̉����X��B��iWtum�\��P���PH1i���g�=�-���o�b��	��'��6��.a$2S
�����}J�n�o E�C�=��]kإ�7�{��G�L13^U8e��U1��\� �V�7J,���V*矙�2�[�IZ0�UY�岖T��}�t� Ut���]��Oo>fjX�y��I�|<G�#�+
�����H�lj�1�{��P���輫�jB�`
����U]�Ȼ��5}$�U�/������ϕC�׭��-����IA�>?Ǵ8z4�$�G� �j�j��uFvn��͌
��8��2�fP�&C��6E+����W�1������%Ǭ1�����@G%w�`��Q���c|�
�+/?���� )��r�ϣ��C><�m"M�&���C�? ��<����8^|�Y���Z�`7�/N��x��5*W��4#�VN��$(�\��U��4�^���#�ӭ��8����\��_��5��D�jU�e$"�9�;ˆSR�l�8uqBg�"9�4�s�����~��u��a�[������X�z��I�yi2�j-V�D��C��N8�p<'u���;\a�H0w����Cf�g�zn��2�:�tu���>ٔu����o�����n����/ĪsÆu�����g���{�O�7�3��B��N�l�p0�#;�|N��#*��GX��<ش�3���A�ֶ&������E��D�x�]F1=��<�>��4�ő-�d�?~\���_�n�7����q�-ע��r�z���i���s.�w1��k_L?S�Lǈ֘���֟H���O�VP�ܚ����?>x�=\t�e�]>������5���'�45|��B;Ok��G߅������λ0���%���XT$�U�hTdg�&n��$'4�ԭ�UR܉Re�K��2ya!g�I(�ק
�P����\v˜�+U��&)�T��Ԭh8&:apYp����W8,�ča?lf��$��4
	y���!T�uW�
+ۍ?�sz�1a�'��RZID�Uձ�9���䇱�A�j���S�b�C����;E����
5q9~�v�@Ԋ���:B^#�~i�vUFt����H	�<>��Z����u�M)�@��R�*08c����#�����L�rn�[]�˪��w>'ez7����(W,i�y�H�nmo�I�Ĉ�~�|ωv	�M�-�r�9S�c_�4|��l"X�ma���N���OE���GIZ����B4�'�}�V�A�B�MV���r[ǆ�~�1�:�Quc;��u_3-�R��{L4Db�DVh@Dn���1��L�uT\eT\|�T�a��;��	���K��_ĸ�����#���\#=���)����^�����(���1�S��W_zf͚u'ҥ�S��,ʐ�P��P ô	���������{q������;�}M��d�k
��b�C����U��S����"��BH��3�|�5��nTc�pG	���SUF�+xR!��e2�f��gU����zV�&e�Uc����V:	%<��Nk���k��!!�T�#[�H�X�N��câ��)�L`��롛Qx|�=!�U%��te"\
��0H ������w��C�D"އ�[{�~��t�]w������� ��� ��^X���x��O�ګ��x��gO�׾X�d%֮ۄ5������k��_~.�}�1�����-��~H&8����G���}ɬ�p�`pC#3��I�X�Mm(��@"Q��*�y4,\� [��1{�Y��Cw��k�Eۘ����;��%p�O�P�	�w��~��6{gA�Ə��=��9K��ʮ���p�8�1'�����Ο����3܁a+�"�7�A�u�l	�Fi�G��j	Aw��+�$����1�La�̽��k���#�	r!�8�8ذ���g"|*�{ɏ�^�G�KyJ#Q�{�Β�k��B�T�rх5]/^�/6��~q�����&3�D��;���=����.�.�)k��t�x$�fE5A&I\.��A�m����#����_��ǎǉǝ�ϗ/ş} �T+���p�O�ä�3�ؓ�a���ø��'_�շ��@,���+:�T�
��J���Z��e�W#��CM�%����
j��I�iU5K\S�	o3��p�uDT����j��[�M��_��ղ"���y��j��.����*f��#��S����g�]��d�D�E��DJ��\�9�>��Bam䪇(%c\�*#�*>A�P��b;.�m�Z�>!�D�bI�$8���A:2V��HD��)e�+��y.�'����%g+��RE�מ�Xb���
\Ű9��U�*H����a�k�dG�"d� �C8��`��ƫ.Cǘv�s����`�?��D�7���զ�t���x{<�w���6��G֬[�����Z%$�tR��Fs��3�/*JPW�uh�=J����~�^r1Μ{�D|
�Ќ���`!��I`�/d�H�Ƀ�C��CIR���f��dq3�L^��gd������ɾ�71I3����<!��7��<5A"؉����2�ݨ4%��1�p*�B��ٳwG�֭�0�ù2�,��y4<t���3ܲwޚ����G2U� \� �(�]����������c��<��=�8�_~����B�������~�`��<܆���M����j��W�b��?��";�0a"�����@�.w�u':�,Y��~(���78���Ӵ�hmn��쩿>�3~z.�[[$���h8YҾ����@�[�2CBq8I���˯�=��	�>~_ЄP�	��?6v���W^��~;9�H��^X�|>_��CC�,7k�<����O@�aR%9'��^�;~���)E���w?�9�]�AQoA�րp ��������r�)'�ӄ2�X�t!��FL�� e]��3�Jܪ��{���I�%+ N�d�Jq�Y���O͟\"D-[��z>�@Ȣ�P�)ɍ��d2����5/v^�u�c���������H7�2�sw����n]���"�Is`jU��А��N���S������}�c�;b�i3���O�����e�No��;�g�A�}$�H���㤹W#��.�AՓ�CȜj���)5
\rO�������ѫǪ����k#߅�_�4� ��Tdj.K�@H�I�*��B��f"v\���/���d�ڄn��B�U�^�(����~� U�̖����q(��(�� @ԒE���|<���x�LM�s��*q�N��s�j����ʬ����$��<w�,蔗��҄�( I�u�ݠƜ��8�_�P����D DaD�,e�4�)���T�ڸ���s.J�P�a���P�9�O,�*h���2"�_w9(��0yLv�Ԇ՟*�E�X3��]�b�?t=7��}�lǭQ�u��(���1�S}��wn��˯�qBg#�S�@t[�N/t�Ŭ`@^�^�O��t���B��3��)�x�1,�l�*�܍��r:��np�"b�S�xa!r��󐅙��]�t!�����X��O(� ���{����.����b�֋:��U�D�*Ʀ��S��'�c_'�p0���>ف���gӲ�`��]\&]�N;̈́�c�sl�z�x��H�ओ�L�)�0�0�H[;���S|�z�Y6$U���N��ɂg�8�C|^$�6��;���qqճ˺8��.��h���&޸nZ0r�Xl���H�[$���܆9{�iS�"�b�����r9����{���=����ş��g�s�Y�w���u���5|�\��w��j{A-J�zz���o����A�TA2�@�����n���	o���|����cŊ�8���	5ᬳ�����y��K.���;��=��9��@��E�|\yѹ8��#��ᓥ+q��'����Ɠ����h�˃8
k6'�m���l%�QQ08��d�r��Jit��붑���@,T=��5?�|:o8"$F�� w�ހ��s�$^��(�Ӣ�t�3a���&�{�ڄ.�'��"t����jłH�ѣPAvJ�.���W�u"_��X1��$���|m����D�;��Q�ǜ����/�$�W_z�F�c֬����o���C ��\)�x��s�����U�1{w��Vc�o�E����L�S���
�Y���?��|O��8�-�hTla�t�W���&}�v�.�Ra��D��}tzX�̚�CBcA�&�-*"���k�.F.�	bA���6hv�ƀ)�n���*6�� �p�ؚS�/��'(HIdn���et�W��LE�r�\,:(�>�ξ(2G%?Ӹb�W�$�q=A���;����#�/�K�	H<��M��WV���W<��CYD�-�3���N���P6/:�&�ke�� ǝ���x vEC���
OKK6��5��bp{yp۰JI��Y�i��j�1lW��V�����g�`B��f�O;l{���ߩ��x�'�V|��6�����h�3�KD�%�"��FDFvQ��.*�=�L��#��bN	V�~��*mH�d����)���"��F��E�lJ�3����tk�y<��4wQ��:�W�|��{��5������-���O�����ǎ�H�d��Ɔ�<������ҫ��9z�!���ȰQ�L�j�W�p�2sXE�;�bݚ�nلg_x��J,]�R4�U�xC.�Q!k���z�U��J㦫/�y?�1z{���XE�Z)����H&|<�? $�����^��Ƙ8�Qz��'}X�t:G�V���0����[q���[{�����q�%�p��M+����9�~�?��05A`���!��|ǨH$Sb���S�@f�ra�%�1
�hP~��}�����mbM{�W������i;ɤ�ώ�{`0�)'��k~��gL�X�_��;�g�s6���o�M�
����ĕ�߁��`��;�'�������)�r�Ut�
�|	M-M�ʶ���c��~�	~,W�ƻ�t�]u)%�I:S&0<��Ax|� Nc��S(�jK'��X�w�4� J#�|�d�}����X���O���L������ Q���lF���td��1&����.��.��??�l���;�ƊO�G��k�=�~U$yp�n�#kFOo?�<����\��{�p�F�:�![�Q��Gs�Ζ�:��d�4')-��5�cZ���O�+� 9�y�j��7~~e��&8k	)�dE�塞��4�4 !�dE��KK�o4j��s�'Xy�0LN��G�lӧ�S0�
�uI-���P��-�Rڲ	F��p��x����(�=5崓���B��FQ*9ȧ�0m�Ɋa���e�8��}p ��3�Z�I�A�R��p0D&�!Ny6�o>��y*D4I���e.��Q̳��`�*��!�H%�b6��E�mUOXl��F	i^�F����j�ʘ����0t�t��f8�|��5��|�A��WscNC#�>�`���_�=;n�b�=�;UЗ-���� !���^!ΰ�eA�$��z8��	xH�Ш�]J��펛�}L�a��/�^��"�444�w6�GM��0�bN��9������E[T4b)���{�Ù��U�o��h,4�3�Ϲ�hHG^c��'���f�?�Ot�5�����:]0�L��6mX�������"T��\K�A�?�hIr���W�o֣���[�����?*��r�_!
P���%W	�u#�9�@l�ԅ��!��y�p"Z�q�����ͯ~�h�z�u��/�?��w����g��Ó�!'�W_�/��~{�#9�w�q�X���������O �q'a(�@6�.��<�b-��d�s����G�C�{�T�~�(.�{f ,��S,_����r\���hk��v��~�&mm�U�IN>�'i�G�A*1�+/�Xv�HϿ�2���&�}�=8�̳0rT��Ba|��Kp�ᛰ'�%��S�F'+��(*vV���1�57�Q�[�`�Q�P� *    IDAT��!Nc���j���L��h�ݦ�����H��H]VʫD�^u�wz��iqЪO�r?qJ�_������0k�Z%�)G���U/��DOj?+���Y
:	��XE1�!?�ҽ�fV��B/���w��æ�ah�)���B
^'!�ĲK�$j��z�ho%N�_��3܆"4x�!�À�+ԯyQ�e������|��5SH�d�9 ����p%�j�:�������PH!�������tQHa�Ǫ�%S2���mjnD&޷��6��`sZ!s=���Š�����K�U�r��&rW��V���J����'@>I^�,����L:.g�C����r�,"M�HgS�SA����K�?�E&�F�A&���K[:Y��k�\I�yC��!Ad��ɀ�����*��쒁�p�QEc�Fa.����B���c�.����ed���)������N�`8ٯX�$��M�(����͝ʕ��A�����FO���ϋ��@;n��X���]mAO��(���1�S}ɧ���l���X�^�Mqb�H�ؼ�'�rȓ�,GE�Hh�X��T;}ǩr�s*$7�2<R����H«
.a�z!eq�a.8dh�Ys���m4��?��HÕ_���i	�>�{�[q֙��/���U/��ś:O#%���b,z䒍����6�ǧ|w�v3ƍ��f�c�tmꕼf�D2���o�:b�X���V�Z��A�+^��1�u
���<�2b�=�'L�8]�7)C0(0�8a��λX��k�|�M���?�!�)�����t�,��٦��:���_*Fo&�o�^��8�=b��8�/fAt�c�n9Rޟ�n�Q�t4�h�0����Kq�5W�gJon>G5����766#�I㊋�a��ɲ>�'q�A�bS�i>�?�x̟?_��9=R'��C���y���o�}p���#�Rid�d
�|m#G��3ϔU�E��(\e�v?�����D���&�M\�z��'��L�F>��23��)���R������D�H�ձ��!D�����	L��<�UCV#~����h	�_̅��I~�P��qBַ"���t�/�A�K��h������՛�m�ty���]7I̲��?_Х�I�ax�>��O�%r�����"��
�':
�~XLA�6c0U��ߌd��;�`��8�l��*�^2Ŭ��u��Mo���6�(e?�wUHU�n�J'�$� �b`�S�4&��.�"�$��3h�L�J�:%f�K�i�|��N)m���\�D�;��\���2$I��L2��A�xP���#�n6t�U6�,Å\1�h�/(�.��� zF@Sd_G����ۚÆ�D�:��Th�j��G �]%bāJ�Y�&�eiP.�<�x�:��"�MSG������W��
$��� F@݂��oϾw�<��r$
�c��.�V��iF�ߟ�:{��xC^�'��Om�4�h�Nr3�Hf0bb̋k�;
}v{`�(�kWu`�}�
���>9��5�_�x1>��c��$�#i@"��3]�T�$�6�|V٤��&;ª�~>�أ���t�B��j�C�!��*d3�s��)�^�럫z!m3���e��������*>�zC���cԍ�\��Bt��f�4����V�}��d���o,r�Y�3ea�[L����}��fΚ������A�'�x�lM����f�Y����0�/])��7�b(W�+�#A��Y� +����0^}�q�5F�e�ը���s��ن���'���ܹ�����}`A�����ʕ�7on���d]r��9���ufYg3)|���21����N��ܹs��J�� 0@Ͽ[{�?t��C���x�=ݸ��p����l޼I�r �.�׭������O��k��;�#��9眃g�yZ���O?�~$�9�1�Ѫ�$�1��,���?P��F`���}�c�w"��� �:$�\#Qم:�
���YX���,���):��4��R,��2l!%���d�<��w�?����ݴ�=y	I�c���<
F���,�Lz�׺M6y3�t�wם?ڪ�d�>�Z���l۶���1N���%��8�lx��؝��+�����ԡ�����2|�5Z+�P��R�d�E��q:���Q5�@v�Xv�4��"P�F�n"Ǵ`�)l>'7!j�m%����(�e7=�������"�S��,]�yS�P�^*OW@Vt7�5*T(d0iT��˟!PX3��x9T+�T&>�ns�T)(��ĺZ�a���d�sO���Ut�!�B9t��$�(w��.����vӛ��w�D �q0��YAs�.6�|����V2��{��<b�04��6��Y�Uh$2��o3FI�J��ms�%E.�Ǹ[wK3�-�������~��)�V?S,�4"*o�X�@�����0[���_�P�+)z�gPqY����6FE���� G�!�D�pd���[A��Ew1	W(_0��T�5($������1ް����Ή���ǵ���ѿ����o���Ï>�`�ڵX����-S��{[J�A�C��t�b^M���ݞ�I�ˑG.7�m��&�GR�t�.W-*U�����g��
�������R����ehu(���O�|dr��R��u�\A������|-��uI\��?3Q���?��͂��)Z��dI�d �X?Ze�&��]hl¥9�9s:�p��'�O��g_��1�(s��ۂ�_,�.�Y;㵗�t�/�U�Н�t;, !"�x��x����F�����l�b"C�Y�I���y���믓�ς΢�]�5W�'�nX�|==�R@��N:��|?�h!���S�� ���;�~$�5�e-9�e��֛e��5��F�HA��1w�i��R�F��J���I������5�pх?�O<!9���Ě>�̳��[p�7}�<fL�	���/)�w������0~�X|�ŗ��7y�8�r�)�N���e��w�5xiI�F~�L�����a��!��#w���*��C5hr0sbVd4���nZm�#M&'I�Ǵ9��"K�0�X�C�8���O���N��+�k[�Z)Ϛ�o�+�u]zm�^׵���?�I��P�w�u]���n�s���5�SB<.���°5z����cHQަ׺�XW8�̠@��y�|ԧ�h�D(�dX6��Tc���31l��ۏA&����y�G9�A��%[2���s	A����4�na�W�^Ӕ-r�w+�*e� �%WGEM���G��W�+��h�\��j���q�Fz�6HnAE�D��9/�*b��B&�|9�`SXH��\^&~B���� �p�2܁��(��e��c��.1�rW��g�t�i�S�0|"�f��ߏB��ɖ\�}��J\�3�kP���cϦ4��nXy>C�b-m�Hs	�c�V�^/"#۠�&{zჍ�>4i9��AT2��֬�iy3�i��jZ�H�S�����Uҋ��Sp�ND9�U�A+�1���9��A1_NtM=z�
!�?��NM���f�^}q��W���X�?��ą�r�#�$0�E)!�L�u���V)Я��ݦF1����<�p�Nr��)Dj�C��I�����	qu��t۵HJ!mc�Q'��{պ@iI�S�rBS\ ���r7�Ο�������
a Ʌҹ�ݽ�c�]��F8d�de1o��X��3r�aذ~^����R�=�L\ �U�V�d<�; �__���+�,�Cy�_Y>R�ik��ރ�#[��K��N�������W�t��{੧�D4��'�����H'��?������Ⓟ�d2���ke/���+�裏bƌ��y]x��X�h���p�W��C���w�Mn�[n�W^�k��w�,3M�l���O�'�t�|�==[����=��Ja7<~���+�ټ?������~�z�w�YX�b}�	�?�|i(��.ə��_b���8�\pz7m�E�ӧOÈ�V�v�\��.��
��ѝc%*m���8���0yl��[�U�Un�����,�T<Uh�ENh<�B�골�)؄��<�b�&��L��/�k,�.CB6�`C�gy� �\J�J�(�Zg�ZtV�5��3�^��g�8��I؟5��j��F�mT#���?��2r������t��
Oe��jB*=�9D�A13�y�O���Nװ���n�!���� �Br餠�@I�cJ��3),���:' ��"�I�C	�B#}ы�Ԕ�Z0�M�]�u�h�L��ѵVYq� CI�ؐ�M�� �m����J�JB��ʔ���((��+C*6v,n�TA�
����B��U-rxa:ڢ1��C��e��A8`6� �+��)�������%�(�@bp�ۢ���p=���K�d2Y��nD�$�nA��bt[�<R�
<��h�9�5�`�}Hg��#%M��uw��(e1����ZD��R>?�z��6q:R�"V��V�4��}eӏT"������0����ܖʌ��e���y��o[��<���<�����/��*�S�U
��o�H��Pm��aNC������Uw6>��u�{������*�[����/�����Eb�Ah��\,�,�a壯����`i���gr݉'�o��|_���¾�ƜR�z1�YN�*FPZ���VjS#���EҲMX��]>�$p��6W��ԝ���D��w���|�1�?F�g3�<w�|l�l�䷵߬����� �A� ?�`|��L�<]ҍ�|�ić0m�d$�$�J�@���@:�C*�G�<��BT=h�`@�!��&}�.L�a�v��[JY��n�`L"'E����;��@8"�Y�|v��w�z[�����5^n���,G���Ï�SO=�]f�.�;�)��cM����'�#�B݃��><��}8�3�{��7+v�D">,�D8܀���W_z���f�����p�r�,_�\����3&c�ݷߑ2ʜw��(��@�ګ~��Р�]|�!h���>���S���YG�����q��� dO��X�,�������*	�C�4B-ͰVCU�0�ZpSFT�Jp��:���'����r����j0�e�$A��"�?��)�*H����\o5��ѡ�����<��u�s*fvۂ.�4�������SB��Wj��3N=� �������x�ٗ�����<g��4G�T�c}�	\v�o��3�k��	~O]t[#��[q���Ȯ�)1*؇��~�a\z��h���y ����CՖɰ��2\!㼔Vg���A9h|C@j1c��a���JMDq��@�0�r�)�V1�<n������Xs�c&|1��u��hr��3t{�V�nqtT�5��J�p �b�LW_|
H��;����28h����-�7᪛�āG�cO8/��&r>?`/�;�hd2��я����w���?��/�t�p�����Ĵ�(.:�(t�Ť���ӵ���ಫ��q{�=g��)����������o����8r�4�=z"z}�=���N:�h�f���G�n�s����շ<�M͘�f��jmG��Z�-�y׸��o���� ��ҹ7v�m��}��������M�p���#�:�8����������A��k����o�c<�	�s'"Ҵ*a�~�VIXQ�kU0)���ʢV �yҤI����e��d+�5f����q����k��
O}z�e��C��h�F�[g�������o�MoPA	�˪9�����:��߷��,$|m���s`��W.'����vK�Q���Ԍɓ�b�ӐN�?:��,CSS��z�"18 �Fצ5��U0=n��gK��,9.����ʭ�W=D��Gu96����<xv�5]V�3�I	���VGF������(2?ڶ����F�_�f�|�yp%��#��/���/K�&#����_^)W\��� �<���g�-Lz±�ԧ����+p�����pB���a��Q���څq�H&S���={���\�L�:��U��g�ɝ߳�~�
Y�1��/���>��<���S1�/`Ξ{�CF6_D�ۡ)�G��|>�FNKa&�w�d?��<x�=�"x�O��N�)bm�`�D�¨8^�2�$A�(�UD���I�����?���İ��E�S}��N%�A����Ӄ��ρP4-ciI*�j�1�Z�
Y�2�+'>��9�o�k�ꬂj�|�V���߳����������V\���q�O�F��,�� �(��K���#���k�¾;�b�k0c�$�q�}w�K���u}�������/��ɍ3�>�>{?�A$2�6��7��E=�ԃ7����|�ǌ�p��o�ī��P�4�&9�	4�1(��6�B�ʣ\u�`4ͩ�$H�C�|��/��*eC���Aѡ�61�̤�V�hy�I����_BqB�����g�M���[0(;t)���'��J)��������9��w?�n��[��9���'턨������w����{y��\}Ņ8���x7<��<��x�L\�\,�̽�&؞&46FQI�ŝ�_�9�X��jt�w��9������S�xݩ���7k��:9����=Ͽ�r���ճ��9�pĴ
�w�%U�u���9uun�	D	fD��"�A�aP��:"�	��9�L�($�Љ�]ݕsݟ�ܾ���[߷�g���r�TWݪ�U���쳃^8�?�>�5k�`����ta��}x�����Yh� �^�$�?�'�5K:���=�����M���^~���7��������w��tNt5F0��	(�E���{��{�%�_>䟪C߲q��m�w�ڿ?~]�AB����	�@��@҄uI0c� ������l͂��hv[,�/��B�u��x�n�x�E��Gе�=^��SX��l��\"��24W,~���\�b�6���6����O�Ƶy����5��p4�M���=^�,N,��!���r?�;.?k���N�:ˬ0�b����ر�U�e��BVw��YJ2�8\�� �vT#B��S�ܦ�\IF1뎛q��eS��˴$��f�g�|��3����� ��(�N�n��:y��gB�$�c���$ݻ�c�ݢ:�U��bNr#?K.v��ǎ+DB�92�P��3�8�")m���R�U/uSEF1�G�^���9%��b�����шʅhm�S>�l.'z�ٌ��B4WW3?�J�C׮�	7!��?�N�G����G#���)�8t)ԋs���gg����wb�}�ũ���TP��'Zuʦ�#I�	�3�]��;�ڋ��2:6�Y���xv��0�K`t8�5�bRb6cmCI�bbX
No�xw�̕� Co�#�9��@��Va�v�?@�h����q�Se�WC��GfGݮmxMֱ�v�mո�3pۤ�pͤ{QQ}�V������e+0m�MX���_{�|�\6v^]��G���� ��B�5ar��w��C�>�U��ŗK�`�˯#�4!��k�r���,T�;�˯���~�����y�|KIOD�~w�j���f���Á���s�v5TRX�7��Tx�/�A�J���A2����ʊ���fA��h��4(ϣ; %h��6P��!��`V�c�:t�P�B^��M6c�,�d�#k�<:���YI#�v������k�ŝ���
bOu ��|���5/,�o��1>{�m�Cb(�զF̙��,������*���F}}�x����m{S���];7�0+7�Ge�a���T���Z�~�E�J:!ls�V\�������J��߰���1��Ͼ�/��&�����}�ٌ߭^��G�k���׿B�E�:�ϝ;�E�r��X����9���g;�Ɯ[P�u�ؑ��I�7�p&��

J7�;��O?�OUЫ��J�����Ν;���u"Y�dk�ūåz�S{K�J6�Q��/.����F~饗�@�2C'�Hf�Y�e�ށkr0�y�zB�⩬Y�������p(ѓt�j����h^���}���h]�F��
��)���D�p����E�d�����ftF�}:��ڊn];b��!��ox�CY�-�    IDAT45�`�Ͽ��cr�l����7���#�7�m�v���k6W6/���D4�Pk#��0�͙-矉xV#��i9��+V`����r�M��رC���Y|���O���ТՉ�����><ϻw��O?�$��+M`���8@���ѡC�'gg>n�85��� ɱ7A26l��Ņ"[S/��nب�p�m0)d�i!�1���RS��R�E�(v�t�S7_�L�͡��tRE_��es���qLx}����f��w��0�FS�(�pT�ތ����'QS��@.��
�|`>�(ª���3[��)�4mT��f������ĢE���5 ��{^�ްk�@��b�K��DTIZƬj�L�^��)nf��5��d�
g9�V#�+�#D��IAoO}rW;9N���u}ıQzTLDâ5�m�@�~��X�%k�ƛGa���X�b�c
>Y�Gȏw��\5�<���t�45�H�_&������V��^zK?x
*�T���œs�`�� ���}�/�v�?�1��X��99�]r�=#����0�w��Z����&z�?�]8�wp�!	�=���"8�R�� I�ʗ��::5���+j�7����d`�(UR�P'rh1��@���0�A����(��iF��I��'��/Lƪﾆ�i��'���ο#�8�o?���/=���	zc�o`U��y k�����(�}��iz{��33��� �x�y4�
`5�0����s�f�6/:��2�l=�@$�aÎǌ�/c��f�s)��X�qrf�*���	�l���x��л x�ݕx�ݕ3z$f�4�@�:�!�S�zVo�J���N�^r�%�����r�J���<���7w����lGi���tz#G4x��S���9��1����p�h���UUUҡ3h���d�r4���,w�kfU]i����Ss��K�r!{�M�bL_damAf�ϋh���?L�ǹ��ؼhsr-�E�ϲS&* Y��V��q�ݫ��ځ������k� �5�枥����u�,脢y_�
e#jĨI"f+�$
���<�[:*B�����91/!����﫝�;{v�E�R���|�R�c��A�`����N���D4�n�~,|�yt�X*0}&��G���u��N���)SԈ�4�->TVT�+�vm=;=������u�&���1]�t�MG(#�%#J�v�h,�{�󟝏��b5��݀�秱��V���ÇJ�ύ7Pt���m;��x��'a�Y�YK5��ǹ���~�|?�0��0S�$7���b��O>�@c��l���d����UW]����'2��3���|[��h���*�f�h;9�>} N=��$�3���vV�w>EF,:���!��ɠ6�a��ۏ����.��(IRVdF\n�V��k!LK�-ZYa���;�,��<����lhU1�%�S��Q��f0#~�'7�ܨ�V	w�濵�V�~<��5V��F�Ĭ[.���
T4��?�zb�_��gm�=����9�q���c��Wq�y�S�vk��V8�:��%���ҥX��c���N|��Z$����$Z�j��{��������g?�Ì�������V��-LH�gS`υ0���$�����a2�pʘK�+��[�XН�>I��ѿ<�E8�Mky���#Iol���>���Q,�X�b�K��T4H#Ug蔱���PW7^D(������s��)��P��V�J��s���	Oξ����yc.A��n�X��5�1u.���נ���ބ⎥�q�3�Z�े��JL�s6b�`��}��`ޭض�wN��ǝ��S�aպ*��m�`d<=�-,^�#>��u�����S"�H'm���F�o�����qa�s�,�������CcE%vlڊqƠ)�y��(t$��nx��*�߼���)��4pf���xc�p���qc�ב�%�r��������ч��
�Ν;KV����0Iq,�t��;���e�����/\�E'n5�U���);Bj�Id⌕�Z�@s!�qh��B�n��>�)�d��)���1ڵb�ը3E^��v�����9�3�Ŧ�]���mV��}�.GSmiU)�fR��A�Q7-�M�e�F�N�ns"��u���z��؏SO;o��g�u|>?�v鍺���Q���g��a����=���#�ǅ���ḓ���E�"���촋�g�&}�@%�=����X$���U�ʦ�-7M�xD
,�6��Y�I��[l����,Da����ߖŚ]��3x�ｰ���<T�Tˆ��6�c޴�ި�����q���Z�MסC�3@�
���n�c��A���~X:sκ� �{�cp���*�k$I&��6,�?_�9f̘���"��.�3Yt9���r����8��Q�#]p������NG���k�"�X����Q���#���6�X��pj���e��Oߊ�"E3p��-��� )/s�8��ؚ�t#�Y�u��V5ѐ�31GJqӣ�ȵ�.��B҅'��ڑk�w�Z���Zl?�u�FP�ֲ��:����.�[�9Ͻ�5����@�����3��C��G�.�/>��z�,�UW=&J�O�㗵��t��q���'�ǆ�[���ǰu�|�l5��=P�o��.��lڈw���<�o�1�yH���Y�!�p�D��<t� �:��:����u� �|
�Ĳ��B&A�^�|�i�F�s�.���X󲠳@G��c�䞡���u��P�ƌq�LB�&<sRУQ5�<�g3C�^�L�5�!�t�^,|�!�eġ�1��I�����?�Ǫ�Vb��7b�����n������8a� �xR�۲y�Bt��Ƣ�Wc��_��碡1��~���������X���(4�?�'=]��ṗ�����rB�Y��e�< ���>�&���k0��>8g`9N?��v`���ݼ�--�|�h�5E0��yx�i0��{e��r���;�����r�]�<o��?T�y���>���S���~'Zcm��O�#��O=�OU����_���,�X��L��,w�WZMp�,b�Q
��é�p��ߛ�p�E	{�.`yy�R�R�EQ�0kF1,:<&�Gw�����X�, jN�j�ⴎ���פ��;^��kݹ��~�a�j�0�����[C4R����cW����du��S����tB?�v�\8�b�8�@��8b� V��̝/,,A.�C2V��)�>l?Њ`
�I�����v���tC�6x��=�����[Nq�����&�2<0ù���.V}I�zrnzȈf@�7�lP%��US�TY\i���`��qN/DÜ��OƓB�c�O"g�D�f5�F��йY$3���+W|��WN]/K��w��'�K�m����~���B�i2ữ�Ƙ1�IL���>��!8�����Řu�Lx���R�`�.����@2�'O�}�7�He�l������漀�bG�i��f;an��N6<v�LL�e�̘��y�//s�7�� n����dR'V��;"�BX]X��q�
+I��a,�nY���)9;���ƩP�L�����=!W��ŔD�M����;z�4`�Ugb����=o-�]�1n���N�ၻoè�
=��`��Cx���x��g0x0���hnl�����m�?DuM/�!p�Ⱦ 'H=��_p3*d0��[�֢WPP<��F|��[X\Hr�O�6�)��ZMp�3�Q`C��\�.��f��)4ֶ�hU%a�^RǈJ�ĝO���i$C)1Ya�9�U��D:n��n2�m�r��;󭡤X���D�h��69%�C�)�O^�����3�@Z��KfJz����q�i���c�ǟb͊W�P�MM�+��[l¥��B�N��3S��y��ob��k�0��xt[a��?z2.{	��0RM��vk�<�����Lñ=�rĐ�%k�x������A1��b��Q�<�D�G�&ג���G�p�%#K ozS���iC�xyΧ0Ԯ����A�ƌ���?Z4��3e�5S����ʵ��d���7�S2
[�흂��������S���j��M�����_}��=\B�o�/5�dJ����uq�aAgAc��L\��Rf�I�N����?y���Dη����0ØnF�d״��;y&>�M���4Y��m������6-%��i�3,l�!������X��U�A?Фj|?�m3�uIb*�~ �z��`F�u�y.z�嗟a��²>��>�����%��l߾ػk7�V

}�Y������g-��x�o��n�!� ����-���}�v��ޅ���m�s���˓σ���Ν%��7'�c�(�=���ч����E�jS��vc��(V��~�g�<GΧӭr*8N��R{RH~��5����0}�4�x���ESu$�2)���
�S�y,I|�H���ǉ\F�L��TUvd���f�"�N"���p"W5��U����iŞ���(�q�p�����$����X��\L7�uUX��
�~�y��n:bp!��!�"����
,�f��ͅ��N�E�M�s^�_n�c���x������C:G �E�A���.�	h�9�]l�tgg�����A�߄��~�?�xOt��^�w]�/A�LH�ZpL��K˰eS��y�=vDB��B4X����B/b�vl;�`c��tB�.�ۿ]6�����o�!��WI!�9V���Q�{�۳����;!���E���8���ˏ`<�X*�'_��xH��Г�ס�A�!͢9��3����X��R�fb�2�99�n�mg�7`��\�X���!ˤ9�0���5��c�X��T��)q]S̖�KA�s��ªK#����j���P5ڒm�ջ�.��{��r�y��P��GY���EY�hl�`�GKS3��y�lM���T��@PF<��xU�4��:���٥��*� ����?��<�\.7v�ُ�h���ܲ��Ϣ�е�c2
����&���~44����/���B�QZ�p��3�|օ�`���ݿ\0���ھ��nҍ�e��i}/?�l�=������(���%�+++�$�	Ý���^��K!�E�I:;:�.�p�j���HA(��X�y�:t鴣�s�)ڌ]sq�+xm~�����\�i�6�W�t��\�y�q��,��`�r��EO��ײ�hw���׫y�3��jF��c�8�9y vl�Mf����]PZ���z6ZZZQq� �ͰZ�Z�N�PI8:����m���Ե�q�)��
��CZ�t2̤j��0h� �y�a�`���X�z��;IW�7��E��ޖ�z$�U���E�-B�|�d��)����1��L��8���]~��aŊ��'U�D\ˣW��|�v�W����ޞ+���ݪ:cI�4(�P&��@�L�0�,p<��_q������r��@n,bbE<�8~����{�)���;pٝ����7�"����6�%�3&���_����1g�����~���p+��y�p �s"9mЛYk�#�ٽ�1�i�m�<��<̘uN5�-�<��ʎA��l=;d���dŰI�Њ��4!��{"�NN	������i����]#�}��ަ���2�`�\& ��E������ð[�0+F�մ��r����c���Ф�9���d&�U4ΦdVňL\'RŌQ��"�z���2#3�)�12�ICgv@g��|��(I�C
H�a0dU��ތ�~z�l���������HD�s��#�p$-�������Vm��scr����.�4�o%�HAg�!;y����v'����6��Emi����P��E�Ga����� u�5�H�%B���l�^�D:�E.���.�
P�P*�b����]N�)��o}<؊<��H��Ļ�`d�
eC�5���!�JÕW ���@<62�2�\vbT80�L����w#�#��aHg'�V�N������~�?ty酧��rF�s�oڂu&�r�m�aH�i~�0��u������
:��'�?:\YYY�s�n)�~��.s=�o9e�~���p'Kr�6����:��ٙi��g�n����]K;�kP�YY@�n��7�U��t3$����1#���\��̿�5j �1�q��Κ����Q[#���y\�V.��P�В�8��l7�׫7	�0|�I��:��N���_���� CO��F�.�tB�;�oƾ��E�T\��xL5�!L��5�g�h�u!m6��,� �IB��x ��zL��f<�������}�܋��#��\6�`���G�J��#H�$���ge�+v�m-� R�CV��6+<�|�ү��z��pfͺ�>�����Q]��g���p�N�җ�Auu%���j�dea�+7x���Q�X+�m3�!:��'@+J~���I+�m�H�T#7K�d��� ���L���7݄��/Ǵ���h���@ mF���5��XRi�1Ն{n�
#���	'"c�`ǡL{�1Du�yЙ�}*��XE�3^z�^�y����b�~e-��,�b�t�l03=�L,!����[�];�n��avx%},�q���Gd��p�/5�o+|9��X��=ܩi�y�V �r��tzXx��(1q1(F�,SÅ������.�߅s6:XJत4׈����)�4'I2���Pu�x+(�4|�<��&��%�
�\�%�w���→�"�#łU��aL`?�t4��аH%�2�<�TC����n��z�m#����D(+ѨEE.�VGⒻ��N�AZ���V$r� 1�������n�|���Ag�l���V!����	m��%��1usf���Y�+1�,�mF��������{LV�cY�B�(,c�)G<�nQmH�:�z�qA\:2)�9��4�|DUZc��N����`` R4-ț�Y�r1�X��|o�G�����mܤ�Mcp'�5�j���>�Ϻ��?ܡ?1��#�?��U;vc]50���c�Bl|��+�����0����W�UTUU��_��v�AYYG��t�"O6�J*�,Lb҈d��lQ�Ҙ�Eȝd2��e��S�y��\��}��{�P�{Ӵ�Z"25�!��i��l<�6S�]Z�r4Y����fW	u�N#ҩLVu����s����?��X�����Ñ_���=z�{��1��ѱ���8,f���B� $A�N��H�����8Xy9�U��}f	��*YY�Mz�
���#���'��d��_�'��Pk����7�E<�����x�ur���
�nu��ٷ�p%$����V���<{$L;>�|9&]w#���,|�L�:��Y"c-���cmE��!�eg�x��p��q��O�Լ'�ܒa�ŝ]������bv4Y�,FjQb1�8�b�۩ӱR���f(H��KI��;�D��
���0��QUY�{�������L�њ� �脘ы�B�$"L9�2�Hp3���Ø٬MqqX���QBF詭u��3�S��<+z��X��Âք>G>72
KfYګ�͈6���ƌ��w{-��`�g˱��	��2�=b%K�#YsQ�s[�H����d����&+Qq&`QBH�W2-�zZ���N<"Id!�tm0r0���0�������ǁH6	�U}6)�6��D�7����T6��
|Bfˤ�"K�#�	'�u"�U_'GL>[��]H�a�&�&rf����z�N��a:G�V�*��Q�H�"�B���X��jWEl�:z�g��q ��#H�B��>�Pk-2�����2��N��zD)wԙaT�2E�dB8�D<�d�b@*a@,��K[��Y#r)N�#� ND1���Ds��p��㏆۠$�p�M�FZ��Z�s �qS$*�+7���t��o�b�!К��AɣQ�᳜��bpR�a*@2F�+)X��pX��ln����,�1�Xo�w��X��,����~D�1��5�s����3`��p�ԾE�_r���4    IDAT�%��P�����c���yɘ~o/��S���1G`��ޓ��i�=�����������ٳ���-[e�ă��������Y%-�����YL�I=��8?����E��t��}�cs񑂩�3l!d�[�
Q���M�х���\kׄ��uK�d��B������1�дl�����hsw>7�+�:�<'K�����w����L�^=1i�5:|8�y��]�
7���y�"�ٲq���^/�m�Aq�E�h�&�u�A쫨EK[T4�da�yx���n��$�IG�e�st�T�+ƍ�ү��S�?�t��x�tJ�O�����������/q���Kʐ�'��\��E�Q+*-A[0�DR��fޏ�O�G/3�$�s2.pٸ!�K�S���ఠ��a�[�}f�	��0�|��[x���8���8\]�n�:#J�"�=���U�9���YxC}�w��Ӄ{�a<iݎ�(�W�nݡ��p��q���xTT�`�wa�oQ\P�ъd֌HΊ��-)�����N��Q(�f�2��	H)a,x���u2N1
�}�I�]<�uz3�W�W�R0���K���~�qh�V�>��u�$�>�	��=�eO'`�`����ʐ6�k���ܷ3F�=�����Z��umйݢ`'n�{� k����(�2"���,�zER��ޗ���q��g��9L0%��57`�E��q��q�T|��
���2���� �d�)�+�5����a�G0��;Q�,v�p+p�3ap�h�h&�����!�f,Fra	sQ"mpY��>i$�)+��Q��{�0���szE��3��N#�O!ؒ���UT�*��b�C.� �l,�<_2t�D?�����ѡ�#㯆� 6lۇ_w�Y�]X�f��pB/=	4��e���_���6X�fd����[�1��Pfw>B�F{a4萎%�[j���s �
���]�AAI�΂��Z��Dm=,v�A��&�j�WbB<	����e�`�脁иQ��8�ND�����#��B�6�ɀi�&���
|�l��|ؽEH�tr���Z��2D`P2�����Sb�����pJ�z���-u�^�c�u������ڥ�V��������E��_��ǘð&Zo*�+��?��?aA�l[uuu�m۶��X$�P���%"�`T�;#�-UX踈��.�ϼ<�ʘi�t�R���`�����dF$q�Q���6�����9������J�5U��i�2�\\#���ڦA#�i�(��:s���:}ڏ2�D���=��~�D":t�(	e�s�¾��S�?f4zv�H[+͍�A�y<׷����כP��˾á�:8<~5gZ6�ɲ3'�X
���Π�D0v܏?�ĉ�65Ⓩ>įkAkK��x����466���ǢG�^G<��}�� ���k����L��ݧ?���fw�Ix��Wq�=��gBD��uAA��1oC(k�T��9�nD`���C���X���:t�Z�%>[����OԘK���9XY+�d~oB�V���/�w�~U�!�3䗠��Lv���o޶�<�(vn�.�w�ޘ�V�2z�=�2?g|jK����QA����u
ƞ7��wy`5���_���"euI�I6�ͨ1_ڔj��}��`�M�4v*�c:�9�+b�Ϸ���� v7Rt�3*�}�{�]�����M�]���������]�6�O�~_�.��0ݍ�=n���&��bӉ��h/@��j�`5�P(��C��C��N�F��h�D�B�^p��:�m�Ź����WL}5��d�B����E಺�4�Ѱc3>=ǔ���5Z�-��/W��5��3f��솴ɂ��D/ 9@ƿ�6�JR'�Bv�/>��;�����c���z��E�u��$��Y�k2�� Ǡ���&��֛,0�d�R���0X�Cʭxv��P��I�DK���l�!�x�-;#�"*a���B��'�)��F���8.�rIC�L5�ұgc��a���wX�j3l�e�bpY�p+F�V����������E���;o,��N��w��Ufå���ژ	v�O�7�9�\���&�&�펅�Ak�O͛��mW��q(�R�n��vG"G.�s��BW�\:��v�\z��o�w�va[m?V�a..�ɡ T_[$��e�x�3��?���ūѡ�������7߃�=:�m��Ǎ����C�����+��>����n��~y�{g<|��f��%[//�w���=��q����uM�'�ر7n��0�M$ ed��/8����4�8u5^��ٳ'6l� >�snW��*3��b�y�뚾���n��j��GH=��s�nh���W{���y�i�5�!�	��9�:��mc!3v	`I�BB�7'��o��A�����|BX#��˯���h���ۅ}{v��'����h��zt��p����!*k�QP��PF�M� ����FJM�@&.9�aP�]��'\~)n��&���?�W_~!�����v�:�����o�m�����b�z�*<X`�^=����W����>�2�}�y����Ul�2�lZ��4j����"�"�찉��	�:Elt�#�m���ƿL������'�s9�m�t��	�t톊�J��5��I�Z��G����o��@}K>X�N:ɤ\||��q�,|�y��y�#hz��o��:�_��ԇS���'�`�}wb��]��0a��]�W�^R�39+�� ��d��K�b�}1a�<��\���\�;Rrҙ����������<9~���l@�N��R*�!}�c�Cg!XT�k��k��;PL ��]��e�e&A�B�IF��x�"烁��@��C$	r�m�^���X����(H��e����1񒉰؍H��Ŧ��x��x����y;01V�"r(%g�1G��^lX���}|��}X�&�?�$̜=�M�fW9�nb&�51�:aJ��g��Dø�K�o
���f�ߡqSƎйJ$�6��T`�΂.^
�\ 52UMH��0H���T�;Yn�k�kL��~�E��c�>�۲	�-�8c��4�<��6�{�S�{�@} ���΄x����p�Â�Ecv�m.��T��{c������V�%�a�.�ۅ��9�'��>.И�n����+���s���)�p�us����N6��˪G�z&9sf�q����U|
:�O���E�����20��p2(wZ���q �U��$��$'3��˟���������RR�DvVa�	������K��{�`��g�7U��(���_xMlv;�b��?<����;�sÆ��~۹q����y�@]Ԁn6���r�aK��*�/�ò���������+�]�k���{��0�>B&3�����L�\�N��2Z�����*�J�{�޽e�ΈP=���2��;mGͽ�ֲk��ϓJ�y�T��yb$��=�EC x-�v8_��
þ��1㵮_����Y����{�E)/|N����[%0&��!��,>�k����_(F2.7D))�Օ���t|�QUӀ7�yu��� N�9��1����z��$)=��i!J�5�����6l��{!���r�m�����2����u�Ax�a={�Mx�^�pL�������R#_؝;mN�g����He����lkw�#>�^��Aύ��n�p~V$��^y�̘9�<�$�m]��k���0`� ��X��Wy�Çîm�AK�N��ΝP�X�s�\ $�p$�ş~�_���tF5��By�!0�s̏v�C���R0X�8Pی��I����p3�m��٣N���~��8>�v5�V/�
Uv!?�	�S����s�/?u���i�mwN����x��7��H��.y�J�c���k�Ï��-C��FCq�~�;uC��AS4���0�� �˴^���$U&i��1X�vX4 J�����"*&�d��δ!�V�ɗ^�+.<?~�6s�t�?����|�ݐ�U(�L�C4��Û��o��o��8ph��,��ѵ_)ιd�����8Ga!��Ix�N(�4r��ø��ј5e�nm�ő���p׼w�8Ĵ��,�$�q4Dٚ���"N�⤧��N��0*U�Z�����jr�҂W��d��ƈ�Ga��}X�~5vo�����XӀ��z��rĲ&�r��j1��"<v���U�7���.g.z*�ч�>�o�����0rǔN"�P��M�3���K��;1j4Ə)��M7�Gb��bo���#� �t�h�M��ݽ����|ˍ���5�|�Ͽ��V`����Z�9�%k"{8�n����e�aͯضs.��
�o
c��j�Z��H-�t��n�chy	�|p$�y�u��m^|�ilّ��;�߀��Wb���г�&��C��.��K��W�o<�eA�c��n>ٟA��GwK3'��>�8��𨢢._����o��OW�W����۷�޿� V�\)�!%%4#0I�����V�����lCI^cg-s�DT:�~�A

�����k��6Y�5攗�u�Z�����-e���$n��m,�)ΥT�5�Y�58mF��vx}4���쵍���M�E5�����f�Ls*((��Q�t�wF�;R���ַϱ��w��]�;���k�۬(*-���x�QW�O�_��$�0z�y�%Y�s2�d_̅�E�5��O����I�{u��3�<M�v�d�75��)��UiN��ّ�u�f���عk+2�JK
��Ѷ5�e�=u�z��yE�hmkC�]{�	�#�GF)9NDs0�;���!�����O?E^/�j�PW/��Õ8TuJJ���es�w�����"DR)��Ǧ����k�s�<�K��uP��bq	�`����X)�{BQIGx˺`w�jvsR��;T�7��0��Y3�Z�i�)��Vu4Q!�>�D��ʋqB��X��*D�	y6�;���0��"$itc� Ke��&�3C.k.��:ޞ����'c�ʵ�u�~�;�#L�Y�0J"�)i�$[;C���En�fR&"	$Eh��b��jC<��x"c&�^~7.:s0�Jl&IM�oK��﷠.nF�R����&?���`J�`�5�q��kJ�bM!�A��aþ6�\���F"8��A���=�o7 �L>k'�� �1��&��7�A�(�]1����i�̅�C�=�=�G]8��b����Bv�[�s�pE�^|p"ʽ�2e|�b��".8�������ύ�6�y�K; �ԣ�����-��������*8�=���I7�㵡K�.xt�x���0vC2E�݂X}�}*�q����X�l'����g_
�h� �{�Z�(�P�pe��6T�Ż�b`oF����'^��>	�g��M���W+a_�8�(��H*v�9]�&3HT6�ؚ�Y#:`�硥:%��I#`kM#|y1�y�0�#N�M.�Ɍ��V�R��g����6�)u,ī�`���/>��uMx����;q�#w�b빣zO;fԖ�m1}��˸�SwE,�x����d�k�`ޔ�Q��fƑ�SZ�����1�������׭zw��=W>\+.o6�K�[A-0��5C�(����;`HB�d{�۝�3;<��$�i3iMS�t�}4�1���FO<Rgh�Av�T͵N5�д�ڦA$;G�o��,��Y()�i��i2,n4�Yٴ����9�(V��Me�p�T����C?�?6m�(3�M����9��0p ��W�F[$	�����&�HrX<���It�SW� �H���X㌹�0xّfr��� �E�h�v�a�N�I�����P>3����f��9�����r���ّ�G��TF,��z�}��p{�P\\�}�����:�5��~A����([+���m���6��z��p����mN��8�1@���f&a1T&���5��s�~�_��D�C�9S�$��<�NdXNw����W^5Q��o��F8E��Eu֍�@�ڃ�h�4d�oX��7ذ����HY�Hf�a �mF�P�Dh�Q���e����](+.A�h�χ�g����`�9�VH��0Z�Ȧ�P��8��.xn�xd�IX������ѧ��p+t�B$RY�6I�#�F�z"�!����Ͳ�`0:�Κ�5�`�+�`�dٴ*��f�EK��J�)��ޥ�5T����$��l>FXqCo�!���őc
^:���$�nE�ً`�D�m���H;���_��[�m��d30��K�󡥾v�N]�H#�r�-0��PѤ��V;�4RB6dYg�΋Q�ʍb��1�Vе�Y2�C���,�Ȣe�oxd�ո~�HŁ��Jdcj�R�>�8��=�_��w�B$�9�Q�TS�u���'���_v����h�`���Z�5wϼϾ�#^�b,���ԧ�:�kN¯���ܛ�����I�C1#R���'�ǹ7�E��Qb����w��Zu 7]<�]����>�ku�x|�ƫ��a���S�ɚ f=� �.��K�_��h�1�C����6���^q=��TQ��6b�s��^��8U=TI$�$k>�YCஉ]�[G�����׶c�+��ӷbي�x�����uE^4��%v��-/̽1��[���
�}K-6�x7j�]�=`�';Z����@ '�Mx��S���	�-)��Y����������<����wF�1�㱴t���Z4�t���
mFB*�]�f�b��q�{z�Jz	t�3n����)� zI���4����֌f��g�����z6$���[�ڵצ1�5$@#�i�c2�����׬u�\��@un'6�:U�O�22������"�����ѳgo�ړhձc'���O"H������� ���jWC����@���'�2C(�"��l?k{Ԭ�},)Ih��!*�N���A�oΉ��Y�0��E'�;S�u����O�X!~e0[x~U ��d�h�8�F���#c�i�~�b�"kkw��(F��e�Ü�i��j	4`���0���hljBy�NH����U��pm3**��Q֭�7(���Q�ǃ�@ �]�J��TZ�x&���c��9�ԡ��?;�H�s�>�"�=wU7�5kY�.Y�'�\��͋�����)�$Ð����a���㖫�ē�?�ɷM�Mw�@],�'^\����bs�3���}�JZ*q�_��%x�t7�x����/�+���|�����S�ޱ�m�-Ȥ��D[p��0��A�ہ_~��/�a��C�|2!2P$�K�o,����$pr�<�;�r�����j��c/��7��ʜ�9�9:]؜VV]
�`3>u/���7�_�r��^�9�����0ݳb䤨	|՛!n����T^S���)F_r.?��0[�����`�\�BR�1�؏t�*��|z�g�aX���ފ9SG�7��:�ۮ��?N@���V6����%X�v,%E��фU��H�B��;��kw�q���e5�߷�L�/��?�V	��%	��	�栴5c�	�H�B�^BV��o���Jq�٧����1a��>-j�N+���(�����]{ ���%�p(i[�`ʔɢ�8�!�� ����� ��6"nF�7Q�� n��2������
O}�9W)b)�p�,���	�b�p��(s�a�0�ҋ}�9�&^t"��b�AX���5��ś���R��WD{w)z~`��>�dԨ#)l_�������㓡���Y�[m
k3�������zْ�7�<�[Z|��.���ۢ�߼ߟ��o޶����~y���˖-C:�&�e3j�]�Ԭ�,��U���I��؆�mb,�ni���ҕj�j�^\��-��1���V�bE'�B�z�
sj�3��9[�4�G��4��h}�lC���*S�_^��\u/S�n,���æӲA��c1�9��":�t1�I�1l�0a��ܹ�{���F�-�Ձ�=� ����OkQ]�+WT��oO��e&�U��D�����j�BT���Ӥ�CH���(N�B?)    IDATf�L*<��P����@�n���bDZp`�DC-�ٍ��t(��U5A���7��@<E�k�XЍH������\Ym2���M��H�:�j����ϐ��ї���W]�sn��.sV��(/p��f`��c�ϫ�t�l&)!#F��Q�����9��N�e����7=��KO��LI�Ŏ�Pv�y��H&�(.𡩾�:#��spX,����0��iX�v+��?�������w���>�rO1�����nv�i3r�F\4�n�z,���
�����p�\7}:��^zVW��$�	��F8lHDc�7���^]��ݷp�Y��ۯ�Ç����+�쁩�ioi,B���g�}*�l�
�d+�<�7��4ǟX��5�Mw/@S�~
f��\F&ܰ�Ӽf,����í7݀�މ?��w4�]r�ZBH� ��E��Y���� 	"V e�8&\|6��M�+�܇�#a�#C6���vN*,V4�ƩC��5���Eo,ĭ׎�!�BSR��'< G��Hd�Vc�o?	�����FB������M���RR��5&I���Z��P�HFBw�}@����"���z�N��Й��'��Eg��
���it,-C�M'^
��a(Ji�O�VB�)�l�ԦK(�_�?���/��--H�Cp(a8"U��b)��[�,��t� O�P ���&�7T���A:�b��ס�����mΖ�#��5����dSu{�u'a4���!�5�U���$��%n���Q��2�Qd�#��=��J�dZ�J��A��Q�0Ҷ[��LSԔl9��,:�'���uV�Y�p�1����8��Ț�����e���V�s�(��}ۧ�t��H�+����-[6Mظi���X�|����U�Q��!w��XdD��C�<�Y\MsNʂ����o�m׮�Z���i.rR�������dH���k��zN�ֵ9�v,-�E��5}������\�6�L۳���{�9i�J轃 BA��AQ�\T�\A:"  ��ZH$��ޓS�L�{��������ϫ�{�=k�I���֧H�H.�a%�z�PG���C�����=v��0�p4�$�n�ǀ�[J��sE��F���2m&�._��x&9��>X����D4+L�t�"�ݜu|�sp���b?�h�aw�QҩoN��%_I�5�D�C��Ɛ��?��+��5�a�x�vL�>Sf�²�6������A�ʦN��7��͢���' ����S��
����� ��=Ɗ0�����V`�΋�B	(iht+8rN/��7���Ŧ��"�NH�D���G��g��}��f���3Y�J��#��w���������B~�a�6"�j:�Y��(��p��.���B��5~��g!�х�n�%Lot����X��p���9͸㦫��c�p�)���?<�9G������_߇X�td)�I��� ��;�b��-�ۻ���́����k�,���K@����,�c�z�J 1��(��ۆ��s�̀�`�k�آ�H ��;PsՐ�� �_�[�C
.9�8,<�/-����B���n_	��*-�P1JP��L�(@59�S���>s���w܅�{����y$�~6閅lN�A?r�4&�GqД�vq��<��8����k��!g}��^�S�M�I�S<�8����i���hnC�!�����U;��L#hv���/ ��12���0z'��A��Ӧa_&�{�A��AhS��6�����R�$�%Pɧ�ߴ��4�o�L�ڰ�,و����a����9�faYr�$2�A4Fܘ��̙Ѝ�Spϋobݮ8�����|P��@!��P�ȏ��1{F�?`&�Xn���m�I=��ӀZ��V)���}�x>��`z�x2�P����ᵕPb�RXz��i�>qt�"�F��)�t&va�q��웯C5 ��ą����*l��ΐj-�8$�>w 6'�9*r_����C�t�'���������?��\4�W��6���$��c?u	}�G�N�p���t��LQ�H^����ҡ[`'�'�z�\�S���Q�X���#���0`��Ʉ^�����N�>���1�J}|�[7Mc����װ�j�6�>ʯ'�z7if~�
�IE�O����Yf4|�O�������=?%I���u ��c߾#M�>�@��p�R��l
(��ˣ�B�3��kܗ҄���c��)�Z��:u��Ti>A	�1+��X���DU�<U�������nL�Ԏ7݋�W��#�߅��.�����`���۫����25?l�T���2� F{��w��`9ì)d��U_�:%�[���ޓ׍�N��q&ϼj����W��Y�����G!���y;�o/�B��K�|q�7`w��pO�EPV!��X?ObjB	Q�)�����+����.��fM��n�Fz�&4���Pd���l��G���=8�M�TK�{v�#�e�[Ia��!|���#5�PF�Q�`��Oaٺ0�I�MG�^E�����g�^��2��1K!��}�j��ƛx~�(�v����Mmn�=~��8���8���y}'V�Z�W��HZ�桻��y]�R��K,D�J
_8�`\��b�O�P�K���͋����@��E�F�&NyJ�B@>53�������(n�ۀ�����sh�T��+��:��↽l"�y#��<.[x�r
O>�G}�јu�q�����IB��{�C-{},�XЏ��[x���z7
ŧ@�Z&<��Tm۹���M������9=�%?i<݀'�H����=Ԋ��+�'�[�� ���o�`bc�'L���Agg㦆�����-��?�*"�.�@���މl|&u�1eb�]0WDt:���6T.��#�<@Ѩ0�/�|6�}�ӣ�n��oB;�Θ���&����x/�ů����u5�
������Z��!�'c����݄�iM���G�?��un�����@-�QIġgw"�`~�̛1;�0iJ+�Q��7���wQtx�Ԩ���0U8M�.�TB��n���z\��
(hd((>TM/�;��\nJ�!�����o��]����"���I��y�O]B_��ÃW��`i2��=�.X��E���	�\.�����y2� E�;t��W�Xa9q}��iP .I�k��������Y?|E&�@�z���Ի�:ל�#��XW_����3y[]e���U�����|��V/�T7
\�ڄT�L�D�s|��ADZ1y��X�r-�i�?#2b/Tj��-�R�U,�9.)&�Rܨ٬q���M��^r�Ύ�Op�S����% �m�n�Um�'Χ�1q\+���U�`�kطk��D�&�Bg�d�'
��O�!g��hs�p���^�A�]�"���X�����(e��c��~ Ϳ��YH�FmnE�u�`*�s�=��ۋ�~v9^z�1�{����0S�M�b���zn>�5
{��7 �o�+�޺��}�@U��-��A���I������]2@��F4��wt�t��؅�fG��	��$Y����g�bEF�����TF��V�Xtΰ���U5
����w�L	��bI���,�jfٮ#��D���`k� 6�jpF�Q�m�&�&eL���J@q�#��0R��d��A��&�mP��ˉ�<;+������ ܅��m����x���uE_rJi�_�Q+�8�l"`3�K��3�pDC*����VF��p�4� O��8�e�/�l�bn�ݶe-�@����'����1�ہb�֥.��Ο�u�����t���Ƙ`�d����)��a$�l���wಓ��������(���{|�_�������Y˨����&�c�cδ.tG-�z���y�y�u��2��E�X���A�����}�
�p�9�����`C�8	���#����~�M	UO#T�Y�@-1�mp@{>s�a��7z{��˟D���W���A��1 �?����A��*J��8��#q�����B.p�Gi�{���S�`C���'�DV/�QS��<��rH'�8b��.4Ӈ@�N�������ʸ�/��&1��ANKU��D
^��@M��p3vqǕ���+:�b5ŉ���(���]|�g����^��=��_��O]B_�~���?�`��hBF兼e��:�T�����ܗ��<Ɩ[Q�6����jq���_ǲ�v�X}W�\�zB�������R��u�״�׺5j=�ב�wmc��Ov��Q}���?��|}�my`[����'tQ�b�n�H�1��i3p��s"�/8K���h���A�b��"/�x�r�ץ�p�i��@ŝzY�r�!(��Cᐛ��'z�,{_K
�hW).��nhzB`��l߲�ǵK��WT��Q������ng5vU�����b�ё�E��e�)�����;���[C�5��>�,�5������TK,LL�kF�V��rJ�G��ߋ\6%�eǎ4��
F+�]
�Zݕ��zQ�V���`I���P(1�|v7�(�_�{�����f��=l
�Zx!���Լ:�d��	?�LC�Ϯ#l��s��o_q*^xq-n��v|��o��+w��G�C �!v�6�Qh����P�O�sWp��a��epٽ��/�ݿ{w��l�DV�
N�TF�R��BBU,��珞��=�n�V\��K1m�$���E�-Dv4R�,��F8>'ʩ]�7%���:W_~=~z㍘53�\��۰=[E-�.Shy�U5�7�y=��&�yo)�����~E��Ғ��ɯ�F����	0�Q*� DU���d�>�o�j^^�~�Y���ؕ(C�t��F$�S˽�B��
�Y��/+��a\6TmU0{8m.�+Nx�*
�����^��;|�$rX�d)^|{%^z%
E_���h�:G9��n8Q��8�C�7��_��
�T��koa��]��+��w?�_���i(ڽPT�|?Յ�� �9����>��9���7z���_�C?{�TT8���"������-G�����p��2�26lX��/��N8�����[B��6���p�'�jZ	�
�p�gE"8���a�����'7�g�ĝO.E�s*
f��.��X3�w���)��ﻇ� �P/����
.��|��-���Cp6�!�[1��V>8��da�\2�mp�6kBLbtW�Nx�=Q%އ2��R�=^x[��E��q�g4����r��e?u	}۶�&._��Vʄ�><�0�ӡZ<o�*�2b5��d�H�5�Fe��ɓ��V��չ���Jg����ߎ��I�ɔ��z.�zl�.b-�ܖ$g�WO�����qz�c��c�6�ןW�����>u�{��g'N���	D}��Mh�hǸ������l�y�a��al�5 ���$�7,;R��	x���`YG8�����fM0�c�!ۀ݋˩@�0�s�����lC�E�G���lUR�\V�'R��r!�?�p ��l��F��<Y=?Lސ��4�r�&�>��f��U�唂h�}���* �����X�45\^h�*L̈́[uA�Z�3�e|ja!ȶ)X��T%A����f�5���@��̭�.i��
R�D`�Ee�X,�֞�Y��^�s������-�
2�:�	J4��o��@t�%G���(��*l�$��ĝ?�&^z��8���jqṷ�㾧�a�G{���P�Ds�����_Hdq�)pٙ�rkh�x�³�p�q�q�������ptLF~4�B@1���r�.$v�����z��cM8��Ӱm�f�����܎ђU2U��( ��c���8�o2��o7b�̙pWG�_|�?�6�~	��qbAK̄��R�@s(���mx�����o��nX�)�'����9��8��o���&>�)��`ԍ�P��h��=S�w`�����S��S���^�-�h�(6�u˦���0����#,�Wр��P��S�8m~���PM��7\� �=f:r9�ڀ�Ĉ�{.��4����h��A���}�����q����b\���Kx��W0�L�꫾���X�[�{��x�~��P&B^���ő��ᶯ��	������-1�<�\p��X�#�jk ����)��r|+����q����p��w��◗��]�-����	R� �^\�+U)^\�<Bzw�����f�ڮ{��ĉ����{�y�mA�s�P��eS���#B_��#1.��[o/E!׏�]x.~��g�����1�O�j,"|v�r��%���o�sCic'4�)��[5h6,ʐU� z\�Py���J��Xv�������q�T�|�I�w���w�G���xZ�C�����E��'pL�����jN�x�D|S�`���2��w�܃����h����:���f�#�?�%ן[/$���O��>�Z�	�=|�{�Ʉ^�zP����8��ة��daBU��sL����fOe�y�>tO�5Ԍ5[v�b���G�-��=l E4lL�V��g�Z
%c̔���n�=��6v��U%K��T�P�F����5��2�P��by�;�dNq�S|d)�BakQ�d�H*P�α7�N�<'�G�L�5�h�
�c*��/��O��z1(r�
8�T�W� �����2������^e����Ϗ2-E9Ũ�U���#H_�8O%�P�C���T��Dc~�1�fV�z}�&`���B���__�J.��~M
���0��������	 K�Aq���;r�{�8��Cp�w��ξ.�q�刍?�u�X���[�ϗǩ����0Z�ׯ����޶_��e8�����'q���?�،�R��Gdo��C�P�j��t�Z�h+����d^{�q\�ǰfg��5�I ��!@6@.���W^t&���5H��9q�����?-^���I�M��̬	�q.��x�����/����L_��
�q�gq����F6c@�ᰑ2�EscJI
��0��0}R��Zq��c�N�����n���V��M�)�*:��d�й�+N���LL����˲K�5DW�d�/f�7�=�s���NAOĴ���EKW��U�x����6t�Xz�'��3�3��b����5��5��;x����ښ�X7�	��<��C���y�8栙�oj9�^�F�_��;���'/����Ahe�f���Ĭ���`|��� ���Rx���xu�^�`�ȷ�)���r�^��Yőzq`o7��N��������x𹷱����'Eq�\5_��\Č�0;�SzZp�,��'����^X��}�}�"� m^y����.J4��.��VZʓ�t�V�r�h�r#G7ʘ6�����8�M�𦋎|��W�����Α�-+�^1Hհ�_��;wKWE�j����m*����o.��1=uҵ���$��MTZ�677K�����J:c	�kOv��X�����I�ʨ��d���-pe�����1'2�����ǀl�X�Z<V��|��ո��B�XZ�����/t5~Vv���q�P҄�>6��ov�h#�Ŋ������p:�՛w�jm��Dn5�\�)R�|ws/mių{TPD[OZ�R�+�M�iJ�.�q�mMEL���ر��D��z�@ kM�N�G�Ү�"��N���~�w�p��|���ƽ%=��m���N+����ZU,%�� cl���}��B�2>�k��T�ȚD� ����r�h
��.`���]2���"�z�p�*���Sf���]��2%�B�׌&����D��O�L�җrh	:q����[n��� �ձ��s^�/}��0AUS�Ŧ�,�[��JG�jǝ7_�}�4��+(�`���O��Ǟ�h�e+Z�u���ӋѽØ1}
�Nm��%/!�����߻7��gXӟ���y"ۉ���pP�ƅ��n\p�|�p���gu�r�m�o�t|�����+~����1�g-�~/le^S�Z��'7|�:H�0�ۇM;���a�B(h&��F��dء8�1y�    IDATjp��($FqƱ���8[���|�d���Kx��%���	C�C�Y�6��E)��]�|3z� O��elݸ�c�3��u΅�&�pw_�k޺��GbM�8�օ��Pj&���ac���)�ȏ&��{�D4�¸�(��?�v �{T���ķt;�(�8�h�3��0�Uͣ!���1��Xgu;d*v����-�	��񖎾׏j͆B6#�W{���D[̋)�;q�Y8�>$L��k~��Y�ʙ�\�4��!8ʣF+����ލ�S�p�1�Aɍ	��n��ڌ����¥u����^BKHE��¸�f0����f'n��<���6wI��B%���	���������Fq�A�3� �^���ŒW�T�t�$R���f��;��n�^�3�<�%��^U�RC8jB˽]~���d��x�O]BO&��E�^J�/�������v{E����n��n<K7Ǥ��&o<^���ߏ;�h�?/�J�p=�KT̜n
�p�.��ݰ�T���]r��%��4�]�q�n�K�������i��\M~*�*��pq�q�"9!o�Lv��JM(^5�f��*P�dM��=&X5_A>��פ�*�^~���'R�H&˨j~l������`D'�׏|�@1+x�Qx��$��V�,�mpc�Vlp�mۄ�ʤ_֩���l�C��%K�(�R��84脡��m:��|.�
ݥ�
Ei��6�	���in��b)#�yaT�r�F�1��y!R�Ƥ8�S�^6����rD+����l�ۥX�y��X͏Y����	Gs�2:
5⇡�-��GN?J�� NL �W��x�t?s�(�eg[.P��uM��Ȁr\Ϲ;t(D2v�� �r>�bC�OE����rL�5`0����Q0��?�l*�C��yl%t�4B�ۄ�D@\.$
2����皠�b�$\v�U+Ez�����r�������j��蔍%ӁؕP���\6'9�,�L������D(�B&�)�~1ұ;��ڡȋ�@__/�ۚ���aP��~2�t5��SQ#>���~t��0w�~�V5�\�����Ě`s���Z$��Z:�|�nC1�����eK������3���`o��J��p����"�Jh�g��3�a8~P�h��=Z�|;v��(F�l"#S
\%�	d��&�#�܈���<lٺ�Oε�W�~�e4s�nN�T��3 [U���5�������75I���I�B�ZC� �:��5��#�K��BC,��q����-0�*<�:��7�J�L,�\�dKdQ�UD *R0a�d�Z'��w�AyP�5�a��E A>��#��!�A(ի����|C�<���ˡ�r�V��|���⣛Nƅ�J\OKk�-�X�u<���Z���Y�<�t�
����/k3�yr�^� ��֡:Q��,�ɱG�����3���5>u	���G1��݋��a�[���*�R�t3�5�7%�4����+�R��%����f���}�0q|��<*Ǣ��|"�I�]�S�I�������.�3+]$FG���5h:�hn��i�2iD����J���L�`q�mU�Rh��WP0�(�t5���^�Q��� �����`��a��44D�N��܀b.%�;�\+�;v��FzP�w��B���5EdU�.Ӂr>թ�c�!�w��qI�K Z=�Q'��p��a0�#[�-�q�e�Q*���D�;�)�}�(nC�XC��8q�&�@˕�N:5y�p���8���Ι�r.���~�&��k��E��1V�Ř4�Cg1���֎��$ڬ�e�9�px��d{dr�b�@9r_��NFl[Mx��� ;@Ŀ&� �ѺQ#�y�R�^�cb?UNt�y��&:k!�@�W�cTGK�����T�>R��!�;&dD4���P��Ō�P��C�4K���u��V����r��52@�`A�ʒ0��x�p���qy�dL+}��!8U/�,�e1��M�%�ˉW�@��*�
U��ͨ�T�.e�gY�Q��ev��/ E6ǤdT�\��r�?�.IT�TJUl�N�B��Rq$�芜&p��Ǘ�ǣ��E���y04�Dͮ���������ڌ"T��2qZ�6�#�x>8����0m2��񱚁|��|v�"QJeh���PP,���@���YC1�A(�G$B�TA!��=/��,3��ģ���L$�2±�(ە9�;e�B.���E������<��B�Bv����ka���}+E^���`�5��N� Y�/冣�j(�T*���&(���#1�q��J^6iD��^��(�1�)�D,*�vX#�fʹ�*��z*���è�"I��D��Z�+"�����+��6�~
�z؍�`�{����Buxd�K�J��'4<��s��⡍���p�o��2�?���J��ٽg֬^-��T<��Z�Cn:�qݾ�tq�e�]vdsz�@�:��9`�4���;��:�:ۡ�X��CM-�\�n��ArUh�JZ.��RA��i/å8Q��e�� �+�zXT�3�H�G��Qs�e��'�֤�E&�(�0:ĩb�H�6��;��Y�4�`'�b��N���"�>w�\�b�Ѱ��<�Z�`+G'^�`;��1\4Pu���1Y���G���!Gm�B��F��=����]�f�i����:24�v��t�ao���pTTL�b�ipy���&��:G�C�j.T+:"^j�QT��p�4I�,ָ:a b@����9�y&E�>�����Rx�N���������c��E�Z�TB�熮��-�)�ESc��B� ���ر�⸷dz�3�u�h+Ȋ��%�S,�E��o|	<O�c؎1]vM,j�.R��i�:�bv�d�T�+�h��}LytH�㾞;���פ�'��g)�q�/�4sq�BJ�XB��_ng��=3�;l�^K�E�Db� f�Ţ"�>	�w���WAUˉ�o �	T�2Z�ʄuy��Y`PȎv� b�%��*�8�[gA���Af�ت������Z�gQ'z	dH��
?3�;G�'N�\\'Y�Fɑ���	N��5E���g��KϢ�j��R��"�#�9����g2:)�F��>�������2;��^Bk[��dq�Z��Z�E"ӧ)eD�a���(��0�e��VAT.�ۜ>�DƘ�4c�`Uj�$Zr�Y�q43l�1��5(�[Y�!Y�\�X��ү`!���4�,o*�����|c�Nd�C��7�#b
p�(B>3�.N���LpH��ꍖ��<����N�)R+A/�1aB7
Ų�o>��?`�S�S��:c'N�D��i"M�,��2�;E�fG!_���Gc0���=8l����z�%��������ʄ�����������x�u�ڻ
G��'��푛�o>�8
l�y\��I����Ʊ���W,����Dw�,���PԐn��/�kǩ9Kp�-q��jn�9-���#�|�� G�L��g�0ZHC����_�EU�RA*�(^�
f�LDB(n���g������Q2`P[��q�����Ξ֧�L
s���k�����}܃)�G[�x��7�P2U�\A��p�lbLvT0��3�Ko�oM�i�-�=~ٵ���2����#��,�샍��k����)�N���BM��T}(�@���Ά]V}�L!��4�� U��� �5��8��A�uC�;~�D"%]w�Ng�-@%��]L�8��\��,g`���U�P�%�i1���k�gL���ym�6�b�3/c�=r�re��P�]�2����t�~���I7����*�t�ğ�h�#�/;�,�8���;�*E�S�y��G������p�^&����h�����(�Q�^*�����8�~)4��Z&��l�C�����UEm��h2
�'��gW��z��|x��b` gwD� ;8"���m��5���������� ������\� /-&E�D��R��",r�TyQ�՚|KN�8a�x��\�L�c"C��X��e�R]��*��^u/f���RY��z�D~��+�,�4SN�d��r������y<��S��8]T++e9�oG�P@ޓ�z/U��,  BZ����z��7j��Dcs#��;;j�
Qq�7q��9474�돌����Ʉ�\{�#k%��V��q�9�ikm�����k��Y�k֩0٠���2�~�tI+Ѕ�Z�ԏ�He;mB�T8y�Z��r�u�Ц��p9����hP�|� +'\ք��	�q������T1<�6����0�����|�
E/����#��t��s�k�ۙ�C�2�?����z��?���ۋ��c`pP��x�TZ�=IIc@H�G��KPlg.��z�>�t4��M�����g���x3S��b8�Ώ�^���N�(�j�BC	>�u���}(hy�}N�;-]C8�=*ǘ��$��@w9�	E��\"��5ttĂ0��������)3��}�7�f��+إ���޽jZ�;�Av�VU_�̙31a������ڵkk�	�$Q�v �)��.�o����t1�������=^i��o|����[a���_������e}"�j#j>�j�JQ�^�$��M8<Iܷ6<ݲ�����p�142$�f���1�����_
X��r�3q���-ʞ��fjV����Վ#��r1��H�W��SUD=pڌ����7� >Z�=�&��g2Vl؍g�X��J5g��[*U�Hi2�𺹲�I�
�3kR��,�m]&T�<�M2�����+��5�����>�e��n��B�t?�6����&�3��L2�sW�B��a�΄\�P+��7vR�8�
谘ga���F���		W@\T*ex�T�VA�.L�L���8�g�g��dV,�Ƥ�ʰ(�������E�7����KA$���_�E2ϱL]j������c�c�!�E>&)N�8�*��P\�7<��x�c�>����@|L���ǘ��1�E	#1�A.O�����]wҫK!S��]I�-�E���>�Td6ж5��ZN�\���5-�~~�[���!᯳&mm���H|�|�L�ly8��hji���"�9�0�HJ�}^L�l8�4;bS�k���&Y#Ջ�\<�\gr䮺����KU�U�\x�g��6��@�F�>|_
Y�*�$�fup/�M�\�B�ߕ1��6qQU467ax`T�͸�.y���~a�H#S*Iq�8('���űD+^�$yY)�����xb�F�H-�b�ʃq���K��uʑ3'����s����T&t�[~��_/Z���D2��=�.��p��P(P�z<�ZMχ��<���q4y����(�etuw"58��y.�]�S���UG�Z1���X�N��d1%;z'i?�I7t4��/���`���Pv�� ycm�aS}��T�܍�?���?| �W�b4��h2#�TL"�!��EL�2�P]��V��3�yV�
�����+W�Ċ��Î=��v�^TC�X��[�(��5GB���_5�)�v8{���|�����xϻ�_�4�*k�ؗ�Q?(�ń��B{�j�i[p�汣���MS��o��f₣g�(�dbMb�2m�4lݺ˗��_|I�8k׬�8�K?ٹ�V\@�ք���y'��]zG[3����� q�/�c������b�����8��3�u����Qh�	�=�\�ø��ȿ���40s�sI�[;yӎb�,{Y��P,X� �2�T��.�y,����A�瘶��>�TE����l�H��Vy=2@��`bb�t���Ȱ$��;��{�0,�F�iZ|
�@W{'��)�4�7!�Ϣ��E^���cpx�c��y�z	��ry������CGg���3�?Q,���D,� �ص�L�L"^�j]�v+"S��uM͍�;`Q�cʄ-#�1KT�F9i���6y/96���(��FW���mڴ	MMr�x�eW+�B 	J�IմR�"S1RGi1K�\[������K�[%oi�j��~%p�kعy#
�4<�"�UđhZD�ͺ&�Z/��i��'w�.�4wa�Ν�H%�+!�ә���e啩Y,=6%�Y��.�[g��`��������),ĥ��3�\��d�����#���;vnƶm[���h�>���.r�kĆ@�/5߫�p(��1�~�q]ݒ�5��{PT~�civ�Uk N��r=0�[
�\�(�lUy�Uxm_){�"ʓ�ߌç4�����O��I2����&�����G�9n��QVl��#)455զM�fEο�ٸq���8��E�t���)F�p 74*cV��RQ��
��z�h0+pkyxٱ����]±��4��y�:xB>l�)���	*�F�(0Rp ^ґ�RG8#����8pr;f���jC$ćkV���g�y&F����e�Fd��*��,� ����I�����?����rbջ�$�EZ�Pp8��G��/,�-6i��_w)W"��2���WZ��cO��&s>��g�	<���w�)��Vb0�>A3s��.��$U�餡�45��!xC���OŔ��l�s��Ɩf�����w��Ǯ]{�b���572���
��&�e��M��[aȺD�K(E�N7ej��ي��F�f0������I=]��׋ݻ�bӎ~l�O���)(���H�ӄb��h+%0o����H �K��yb��H�ߣH@���@Ώ��k^��$���}�&�k5I\����q*��jU5���C�çZ]?w�M��&F��Y(�$p3�2��)�K�zhޑ�c�z�%�^���+��ʵSc�&�P̏�¹��\��a��DjԢj2"���qXc�:X�4H~'�Ζ��/�H����)���M\w�L��.b�B1(���7m���c�|&L���I��
3�V����5��?�e� [��4��zS��B�bbO�0�./�G>O&��f�Ԋb��W�W��ڌ�O��u��MC�L�Naw�^��:%�O��r�<���Z�A@��!���t������C��a��󉚗U�G>�su`�]v�F��q`��	X8�^��9�	Bb,�u��铤�ٹ��ݝȤG�3�#�I�G�H��
`K{���8E�U���0Y@9Yw��UבNg����9�p�	�`���[f��XA��ɋE�*���RI/	���3/ǒ�F�y4�F>�/>e�珙2%�_�s�]���'����n۶����7p���n{�ȝ@|dݱf�:0ؤsp&3��H	�'���*£%P�'0�ͣ{�AX��$����(&���hE"�ĺ]���P+fe�Y��U�S�9�#a�P��H�frGO�Y�`���a�Tg,�U�>�9�-D ��o��7�~G*���464c�ҥ�2 ��c��@�͎�����W��y�Pj�;�	dl6��g�v�[�S�����T�����V6g���}�����c[�Ϳ��W���p�a�ކ�+*��d�J�}�é�� �Q�V�#h+Ñ��W��������]ѡ���{p�-�Fo�|ȡX��uE2�3Is�.t.v�����[�$A�;�"�`5Q��Q�Jh�h��q=�K<�B���?���������q�%��Q�\�O.Z����FM�B7J��5D=v�{0����](2�i293pr�Āc�ٚ(�c� &�.b�*�KeM|�٢P����W^�tĔH��A����6<G�z.�L�HP�C4��1�����y�8=��fu��*w�y��E��aM?X\��dRƪG�xl��ĀZ.jJ��9�������mȤsr�����Xv����,f�%.�G�����H�CC4*#UN@X�=i8�;<���CO6�olτa��r��_�~�Tp� ǵcϩ	��Q1,Yh*Arܫ��cH����ڃ�{���Fc���ISH#�WTbS:u���n���누��h8蠃0<�[o��H8:�<���k�@���9瞉X^[    IDAT��0��؁����шO&3�wa����w�E
���+\t�e�KA*o��y�gϞ-�ʢ����k�:<�<o�h\y�X�f�CqD#���H| |0�GE�+%nB��w����W_�U����:d��ba޼����X�f�HQ��#�-"�L�y��������c�=2:�t2���>Z��U�VIҗU�Nyi�<Z��w�����R���{����s�d�	9�E,f�4�/,�����W�����7�����h�#�?5|��/�}rɇ��#/�k:��if �����E95�v}]d
�B�*A\x���ޫoa�+1kF��������`�)�A����Ɛ}֏�H;]�l
�J#l�]�����iC�5{#~���	=��&�$�lG:���^Ks֭['#Vvm���Fi�D��5���>D� 1�/�m�֝x���0눓�x�N�Ix�m��
��2���ɢ���Hi�����}��%�7W<�[�7��yJX��m��CS�qN�S��v{.�	�Z٥�R�\rb�8N:j��0V�Z��6`�����Ո'R����w�DÝr"�����F�oh��v�؅C�-[,���NIl�b��w���A:v4L��w���I}��Kq������kV�n�9�[�y4���y�`+W�AG�ݍؽm=��.g�>���	����IW�(���睃�_]v��hҁ�S���e�E��+v2ԏ'��BW�A^x�R�1 ����L�k��.ǈ���~G�1G�TVt�pҩ���޳#i�v;�<l�}�~8H���@H:(&;j7����K.���QD��u�,����{{��4�gdA�x&J^�_���Q��&fI,,~���)k����9�}�b;���I����}[[ۑ �3A[G~��hhj��z!�|H�g��8ٚ:u*N=�T<�����޵cfΚ�L*���~[VU����*0�E�SIٽv��N:	/���ã��$�����|Ŗ�y9�Q�m��ҵ̀��ĸ�V�_�
>��\�5� L�4=�FFF�[ڭaMu�<_��2��]���M�0��W&Q���pđGb�i�����N9�R��@�s}��'�ʫ�7��V���qNUL�(��_"_�[�il�E6�����k������d����*	=��!����q��_�X��s����׍�L/�`!����P5����"�b�N����p�=|�"������8�,\y�U2�ij�`(>���A�|�ɲ#��ǥ[ga������rء�я~$�	Q.1��s�F�EF3q�8�������������M�s�>�:����?,]��W>����Ʊ�F,5 ��r�gS����ْ8�7���qx�{P���x������q�5�V!�e	��Qv�VCV��I^mYG�h���$l�*�p�#P����3���WB������6lܶ�pN<�t鍦R��ʕ+e?ʄĀO4'w��Ӧ���]"G�L�w��{�PD>�F��`��X3�!��A���Z4����`�7��&�\t�wnz��h��o�\�i�������5�j�`s٠5�"��.�:�x����M�T;q��g ���ge��Λ�='O����^���.���$�C�Xd�f�8�|�vr��}w�7��N:�Ì��c��]l��X��iL雌��&A�2`tv�H�T�X�i;�|(�8�x,y�M�⎻�jC?�J;*N/J�"|>7�D��E��DT.�|� ��9�ҁ1a�f�.96���.\�Ï8�_����{�\�ulڴO<�]v&�L��-�l�+.��������t��tX�X%n�u�r�9��k��Lȗa܄���7���Y��	ֺ��������_~�W1�vx�,Jd_|1�O���7~Ϛ���������'N�8b�ʢ��	��8B�0����Hq��cb�d�F������㕗!���PD���$���ᚯ^���!<���� ؑ��g�}^}}	����O�����~����=��W�BWO�lڄ�O=s<���oп�_�pL@���\��U֗�|9��0�}�uhhl�?��}#�Â䶴j(-OЖA��j��&t�chp�LK8�:m?�(���Ǳ~�&���hTeZs��'b���p��`۶m���׃�{�c֬Y8�У��O`����p�Y����'M�ŭ����&@�, :p���<�֯_/�eAF������oW]�)ӧ�[���\��2�N$G0o�<̘~ ~�a�]�n�'�9>�o�D|񋗡��?��Mhhh�v6���Ĥ�����A%6V*���ĥ_�����?��"A��MĎ��Z?�����;o�)ǂ>����'M��#�8���ϡ�x�X��bB�'�uNߥ�����G�����M�sd6mz'�<~�Y�>���^^�m	2DI��UIG6O��((�����ĉ=���0r��8���X�"�I���Y�<+�3�Q���bJ�Լ՚�>т=���#�yƄ��#\�,���hj�I2�Fx&��G�����.F�il۾�-��h\F$qӧO�= ǔ����N��C�r?�rfV1�c����8^\���6T�1T�U�8h܇N5���vᅗ��	���n�ᅥ�oZ�����LY�\f^�eq'J\37ȓm�В�0�'�N����X�E��#\Z�('r뭿�=��#APғ4-��hmi��wߵ��+��7@u:��Ԋ-۶cҤ^��	����D����̼�=�|�m�|x�xw�Jx��?��w��;K?��>��C���K�����zH�bBGFwC�B�c��$���b�����#l1������?�Tw�qz�Q��dr�/�@CgAsLؼx2�fw��#9�����/�g�F��g��1�xᅗпw�t߲ct;%�w�18�ē1��p(`ј`ù�9G^��g���Ȉp�����I8�?>N9�$��y睖��ؘ���/c��}x�G�[�螝9�]�N>�T�p���}{�1k�m#�΃�?A�sz�	�?er�mv�{�gp�R�=��R�$�Y�^��9�ٻ�?����p�EOݨ���g������L������Յ۷c�ܹ�w�Ax��w���U�d����o� B~N;�L�<Ã����d�é�Wv.�y��E�)�f�=+0G��J�mmطg�L���&�����OēO���]�ƀjU��L�g�~:fL����(c�.�m۾Y�~3fc���X��-;�����܄/}�KhmnŽ��/׵`�����:��Ǐ�k�_��-[,ѤrY�9��|�X��ۭՇ` LQo��N�>�<����j���"��A�Ă��Ys��)�� ��& Fp �}�����:����}+ k����������nV���t��� �<�˗��ի�����N�sL����u��&�̹Rv���9��c�?}ތ�4��w>����5k�:���۟Y��߿�>�.�"�O+�t�E�����Fh�J'Mv�/X�;7���]��ʽU�Ĝ��&�l�ꐮ�Xv�d6a_6��C>��H*eD[�`�*��m�u�3��:����v�X#V�Z-�ӣ�9#����b`h�BpR��R������e>�N�T��#q�����|vbh�$��
�=y��(@�Z	 j&0=��<�?������w�����ӫ�IԃP�������/&�ߠ�|�v��U؊C�U���7b�ǠV)������v����x�)99HN #S �)""Ȍ�e���p[m����j�m�X��ޖ,�Պ)ʠ��1	C$��p�ə����n�o���z�������;>1�u����������{{��Sb��&_���7}�<�,V����)���d��v�|}-X���E<�u֮=E<�}��I�"EnxP�'��,|��0����|������֠�5+F��wb�;��\������ОjCP,`n{�c��H�ujb_x���N~����p�����Z/aL�>	��ἆ�.��r�|攼-�<-�E*e1'No��9��hL~���FK6�
g>��[0���˿|UēXx&=��;&.��2,[�\���1Oj%�?��\)�����x��bc3��Q\iN�_�n�xX$Gz�|�X�@�}xx�=��m�.����i��]�f���w��x�|/z�^x������}ُl*)�wȨӕW|@>��o�B���Is�;�p�y�a���xj�f���뒗eΝ�jzk4���˳s�����o��G0d�'�t¢����:��[?,�^|=�̵���� 	��f�l2����y_줰�2��E�Ʉ��ysq������"t��bݩ��ē?���_@f�Hͫ�E��]|	�<�<��G�s��;g��K{�܅S7��)'�K�E���i!zvp+V,������;�G����-��#�8��Đ����>'����fp���`[�n��+�KڏEm����Xzܱ8�u��?��f��aӹi�^��_-z���v;:�ېH��8'x�p�IbL|�{��+;^Bk�E"Ucc�X�p ���bt��A�)����7:<"���ߏ�����JX�h�;���O�+_����:��l8}���n�iɆ&�_�����VB�T��٣��w��ې��Q����axU!�"��J5�4e��Y���޵8�c�HV� W̡F�3���z&�|����R؂�j?�Nd1:�A�I����J'�|TG��3z��>�o	�dA?fredZ:�h���J_}m���J����>����������·���Kfz [�lA߼xfܓ?��^d:�Ş�^l=�G�7��o"�2�kpr��S�w㮸1���z��O��'���J�CՌP���V>�j�X{�-�$��.N�-�b�`�w�"|�#׈����ߐ�իWc��C����M�6Kn�?3C��7(�,��H�l[��'�x"�~�9L�����#��|��=yM<P�Clry,Z�'�t�`{�}��u�\�D�g�غc��"D�nf����M��SV�����~�R������ �8�v�¶m�fۼ!���69���0/H/��X~���7}Xr�<�~��XE��5^�^�g�q�����9=s�f���� F'�%��y�ft�w���$��]p��Ӥ������+��MO햛?,^�O��	v�z�mq�{�y�]q�8�ӥ�[{��1��sW\q%FFG��O`�[����)��{�y�3�:S���Pz�4}8m�zI��`���X�!��I�W^);k$`*�F�ˮ�B��?|��X��`�#�W, �q���Ӱo�^<��G0��;_}M����_~Yjrӓb��yvi�ɟ���F�I%�/���w�M`_?sߌj�9	�Ӏf�+�j~ܑ U9��U+�c�Ȱ|�
����K���?�_�ډl*-�C����sލ���=x��H���{
�������x�����[�K"a���V�^��.�'�����_H�&�͈���y���e�o˖��28d(%���ǯ�j����ۿۢ�[\x6�����5����ó�m�����O_on��z�\y>��tKBR;lW�}s��Ā�����7^ۅ������_��V��׾!{�;wFG���eDa���x�151)r�T����ڈ.�P��~���e��M:��;�m�����5����u%�w؆�;�K�����l'
n�|�@�*��ɩ�x��W�̫_F����^'�����"4a�q:k��.<7�j� �q��¦��8�K��:��>h3P�T-��c8��cq�1-X��'C�V�VКM���]ri9y���$�ɶ�9�se`s��⇆�����)��T�<�ãcxsߐ��?��O0��q�����PnuP�"����N^8��%�k�e���wl�����������7~�ln>F���"�/�JVKӳ�I*��k-� S��c�p�|�����o��Ov���v|����R�	i��ux�:��{^Bg� C��K�H�mۋ�H�"�O^��{�bt�0��իW�,�F��7����K�摃��I���B2��+���-��l_�Z�A�B�=��4-���u��6+x��`F��΋���!���t)�b�ؘD6n<+Ws6v>�:��
!�@�'ٱ�W^�ߕ�a��T$DMC�����sH����pxt;w�C��_l�IU��y�{N8�ģ:ɑ�g�up�Eajz?|�a8tP����	;-��>�h��ý��
~"�R�y�O
����Cw{[F�dh	Y�;�T��p��Y3Et�Yg	Y�h��&���F�7�$;?���s�͝+X𞢇N��?�O
���F�Ù�:�q���`�ҥ��e%4#4�(�t�gK����<+d }�L�x>,X��/�pV�&/d��a��-�"����j���k
��㔔5�ϞCxV�\�##���ş/Z�'�ty�YK[;���(�(��Ƶ�݀�O\-Q���:�JK���0V��֜!^���ψ�Ù�c޼�B���ˤN��u%A��q����cr_�Lz�������'>.��]w�ݬ�l,HT(Na�	ǋ�����+/=/�pG�\>t+V��n�--R�W��a*L��a��|i�����X���'ƕ�F�����S�A�|5�;^Ź�#���?�{���Gj3x�����п���Jt��q��\z�����/|�?m!ܿ<w��߁�{�����_������&1?i"k�(�BL�p�{�C�����JS!RQ��=Vα�05�9�"��+D͈PsR���+'12Պ��Oc�͢���r;�b��/�Զ�FX,�<r W�{��8�hF,ݔm#��򥋱w�	�� ؽ�-�v����[p�{�ő�1i�a,B��6㶓_ڎ�`�Z��l??�zS�ؖ@-�`Tp+c8q^�m�]:���z���~�k������M�&>��X/J�~��N��r�:�B5��{(R���4L�����kq�?�s;��J�=��E_��s�����x�J�ǽr�r�0oz��}��`��\���p<~&/y6-�J9�S׭�C��-����7%�}�g��s��I!x����!�l�H���t�J�űК��,��T�zq?�?�$�����q�����×�N[k���4ãˤ��-nw�}�Ѷ0z�7�|�?S	$e�q�&1_���%\����_��x7uaV�������_��KdR)�l����_r�e8y����Cg������"���I<�ԓ%���Bb����H���wW�\&6u����z���x��'�_��IORS--��K� ��~��<h�Q���~7>,a�C���js�z��K/�B���v��G$au~��Y���><��#9"{�/V�����}8��Ę{���{$�7b���h�����A!�|��^��	ǯ�:��-f���|q�6,����3i�2�N�>� ��@��t2!�{�,��C����X0=q��~X҆��<���X{�:�v�m��׿HT��G���7��(s�ޔb�г��g�õ�������{����Fc�����F���<XH+-�����G>r3�/_�?��ɔB��>�����+��C�0�Z[[��,1'K�rˇ�fͩ��OFe"��6�?�-�w��m���șH�e4����]w�D�n��cHe��Ӎ��Qynي����3�A�;vM�3��яK%�o��;*"E#������g?�����gZ3���;��!��?���'ڶ%���i�!Q�Rh��E�f{@��;�E1��/H�5d1�ũ)��/m��jp[[px2�CLU[04�B-م)�z��N��A�L{�ƽ؅*��ݸn�"|�ҳ`��V����mR<F���a����d�r������
��A`��g?ۄS֬o�y�U'�$�Q&��Ժ���W1$�ֿ ��^���#X��ce���{������_��7�'>��h������̇cs�!m$|���lŷ{ոw2�S    IDAT�0g|>u��8sY�x�p�eW`ނ���K*^=F ��/�o�,̊�ǓҐ.�k�P6��A��y���U�0U��u'��Z�yJ%9؞�^��)�z��X�tP*�m;�<�m;b���ޏ�&""�®��f�jQ/��*K�P�ʸ�ҋ䰣�������ݳ�Y4nHb<$I��X�Cg�������7��lH�Y�
k���%^"c��0Wo6n��#B�%o{a�"���4[%W���S�8���M.],�!bĨC�O=���]n)�����*,Yr�x�ߺ�.9hY��u�%����ò�_�x9���� ��$�˖cbj���%� �k<��%����O�(LG[��ʔ��.\{���HB�;�C�A��	\~٥�=��S��������5��K������7�#�@�.���7vcӦM�=bE��r%��˗ᢋ�/��^��w ��j����?(��l�����=�΋�mK/|��Ǣ��>�NJn�	���/�/���|/�b��O����O΁��n��=p`��W�X3�;ഷȖב�	����{���h�������4��|��_EGG����#1��՚M�>��1"�R��"Z��[��흂�ŕ�t��}=rxH�L?��?ĝw~�|���(�|	޻��֝�'T��������(�-�E*���i�\t���b�+��x�1e�ɛ�g��'?�Ww��?�s���O}�C������i���J��������?�p��0;�cjb]a	%�@���چWq�Bd$ 3!U�~�0�2}�C�]ҮS�ּ���4B��W�p�(��E�(ͱ�݌�����2�睺׾=��
��0�3c������_ǂc�b�i06�Cd9��0o�ݝ��¸��%�,��d?��/��{�
<����ZSH��"�ҍ�#c(�2�n����GCCw~������=�Ǜ_y|�>���J��`ZT<�'�q��c����6��G`�&�(㊍�p���/M���~��G� ��Jg{6�|\���9[�� �P��h�ӻw�q~�^�]�3���F�W���|������x�z���݅�s�q��AT� e����v����(��iz!B�y-i��t��ҁ����H�!r�i�x�B�������GX�d1���j9���ۿ�P"��>��|�\ǜ2S/��p�2�Ӳ���<�x���I`�rU��H��f{[�s��GGư�5���K���o�|N��h���n�I���9�}�C�����i@�������#�~�ɍ7�$Q��~{��-�`��d���l�:�l����G�ʤ�+d�يu�	���B����>��6���lU?�\s�_x�|��_�����Z�D��?��ӱw�۸�{�xn�������'���) )ң�N�"y��/8g��.).cj#�\dZ�P	,�NL#���K��*z���qd�����-�>|� Z�)��!e�96 ��:���k(�ʲo��TЧR���g����`	[
%���315-�
�MO�2�D����7a~����Q*��Q���fZ�?a�������(�$�Ҵ�[��\�0���t�sɰ���Ə~F渹f��)������Ɛ;�h�(�J\��g��(���-FJ.7�Tv���n������g�7��uδf�]%�w؉=e��ھ���P��e�^�Y�M1��	��.�Sȕ*���iD�s�����QM'0�������3[d$)�(�Q�&ng���(���^�!�偩������K�D�Q��8�P����Z�`bj�������KU�޷����p����rݱk��<���?�-��(�Ǥ%+_b�}����Z�c��é�5���������|���&��m����SN��\w����-�h�`!,�܂-`q��%x��!8A�kp�`o�WwW�q�Sק���y����j���J'(X�����I6P�X�
��"`�Kx�,��>��H�y)�,�RǏ?a��[NĤ"_�OW9���5��q���L�Y����a��6wݪ���%��Qݟ�^)c��'�{k݅d�U*y9ݗ�^?l��D�����R�t�w�g�>q�;~"���K]��k��� �:�8�Y�a���ϱ�\Y6{I��ӷ֓g�{��J�>�۰�?:;�(��+���ǰ� +����<}�j�nȫ�6P*JY]���8
�*sv'��Q5$w[�-Y�^f5�>;���vƍ�{dV��1�L\��vm^��o���F9?!�������V�P8�6	�9&z �ڵ�Cþ{b������ۼ�WJ Ć��I-ki��#v��f���2��5�
⑫����K{���ЃU[♾��':�m��}�0����ެ�[���l}�^�7�Ⱥ�ydB��	rf����겔�G�I��%��'Tڟ4�.�H�X%�p�db!�Ë�\�����
��#�����o<9��a�I��^���/�bI��#`]��j}��l�鑡3#�<O���>�����&�#���}�`��4�̙����(4� [~˛؛*G\�l_j�6�����X\��Ϸ�	\��������b���`�A������x�6N@�ޗ�Ϋ�G|�����Ԧ2�g
�z��[��ֵ�ǯJ�ٜSL�����I_�g;}�;v�;k<$�^�?�5z֘h��#���_�|ێ��~�oB]��^v)��yG�\(���b�"�o���Xno3�&j�����q��[sC����K!�v
3�l��Hc5g�ev����9�?|r*�.���kE/���P�z�OB�>z�=��z��-��u5�d}�q�|�s´\�g=z҄�)��b#&��|�̭W2I��B�<�%��eU��C<*�#����tY��������yw"���Y���cD�J6F�aC~ty]��P��R>�N�{<��ϛx�ۓ(*�����G����.��u��#)v'�/�o��*H�=���q+1��`I��3�r=�F�u6Q1��XP�b��.��0`L����?:��>���qJ�;��ܔ��ֹ��v�#��,K�L��m�6{p>�Z�E0��h���]����J�s�a;��'Ǣ-?,.X�����+�k>?j8���48ߋ��0����qW�/�9��x[���|���
˳�J����������{�յv�Ԋs?�q�V�҇v�$8�>b���=x~d��nMm���	?Q������F=Y���+���bo������,�H Z�f���O�'��d(�?(e�*#F� ��7���Nؖw�)�ǲ$��S_y+�go��~Y��}�H��</���*��
����y���Հ֯�I[�K����v$x�v8��?��p���c����P��d����:$7��iYd�Q��&W�rU@_���cZ�I��������e����&�E� wr��ޚ�ۃ��ĕ���Q���*����N�����Y{O'�S��ՕMn.�S�x�3<]�I�uXφZ3���Gӭ��?c�B�
Q�mivE<��v�������q����a��҈"I�m��Q���.l��R�.0$�j���sK�i�T��e�+yr�x�0����N�if��xrJt��,�����D��6ڰ�]���r���=��v��*?I���a��Bchc1��Co	/��EOf健Y�I0MV����߁ i\��Z4��-�#�<��WL��E�d4���v0j����,#���|J2��;�v��sz���ng)���D�N��"^z݂B��\�߫0IɠUw��5^>A��V�;ҿ��J��|��y8����	z-�_6���_t�����{"ۓ�Q�4�J�Y>H�M�?&x@������*i�dM��V>��dJtӻj&�O���U^�h���wd���F��k%�`��[c2����c���sD�I�<o�7d��NѦ���Ҿ�5,x�/�e�f�K&���D��y�f@���p�A�+�D	���ٰ���0��W��� Ģ�7���h@_v���"חL{
=QO��&�Wh̕��{����ŧॣ��T(D��MYLmb�S����&X���h̸��$������̈\���k�gŖۤ�����G�bȎT4¦�x�����掉���a�b��XO�)I��k�+�r��Q��@�YZ�I�c^�V&a.��8On�8��b�h����1�z3�9�E�*פ��/C�[�W���1zf�9t�>��i�h�fC9�Q,��Xy&|nA�}�J"����&B��� :�m��N�&���[���� ,R�.r�|sD�yc�rǧ�i���28�$��IyZs����6Av��3��s�R�-��ȯ_n�'�;f�X�\��y������!5��6�����qc�j�sc� |C�ɟ���ֻ�/��t7M��@c��?~�5��F�8�U���[����C���*L��Y�+��uؗ��Z�4�6�;o^�p��.e���uk	�4���@Su�-Cfe�����
���I�#g�7|�Q���7}���`u���(&���	[���UA8�cg��1���2���g��h�'Ke�m�N�&̈́�Y�C�1x>�����d��fq�D���ʴ�Q�5c/�-%���Z;[5��}���q���O��8)e:��@�	����	?�+B��&K��
�x��hKL�1�1���揫�i����w�/=�R���]��=��.�9�%�Ł��!���4Zzo�� �[w�h���F||>���%��"���Pd�� ��g����p�����?��K�M����	�$4��ϝ}y?N�+�BƳ� 9Peed%�s�
6k��(W���9���93z���~�&F'[&+��ڡ��N�G��)��y�2bPGX�_�����{p�y+_��N�YJ���i.J{Ѝ�HB�T�N'����.[렡��6_�V�����Bܻ�t2����[:(�1�	u��wm��.��	*���� \��_�T�~|��l�����h�����G���B��I|�n���{w��4?5��1)^�3�fǧ�t"G�J2W���4k�
;"6FG�T�:�!g�
�-��Y��h�n/.12���wǛ��G��Z���M���z�]�Z���~�/�s7_��r���'��M����%�?2�f\���h'�{E��C�sp$bZ��r��g��3�2|�?�鱑X�ܭ�=�Engl���Y^98�y9|�S�����n&p�)����)n�}�{FMI!I��*�nLpjMw.��8��KI�	�Ǯ�0"R9E���S#`�"��@ X�P�l�D��/�����R�u)�S��a����t�_z���yTn~q�z !	�U�U���d��f��ej�5��=�e�A���&�'�)p{T�h��.	�1蹯������28A�+=ctC5:gι$�VRQ�xwzǳ�h=n��arXH�s�3��N��/�mP�(>�:��4��\=�Wd�٨�����d��u.�v^�ʙ����s~��ep*y\w��K��ϕՌѬl��_Ѿ�\���+0o����6L�3y�͓�i~M�)u�z�t{�*o����`�͙${��חew��H�?�J	_��5^�)��K�}�ͫ"�x��OFj"�-c2=*,��{]��KJ.nU`�^��^a8�2\��n�n���\ls��N�c��0�z�M�3U̴�Ur��s�x?L��'",�
��^x�MJA�g�u��3k���#.y����K�rU����OsX����=ԭ�>�N"�?!]i�a4��ӛ�Z�̘��fG�W)��	��O��۝�iI�@+��� �2JE)~����kW���	���
�?��ֺN?���z>����8�-%�� I�G(�l�3��cO�B7�;K<,�`2M��uh�R,�a���;�e�S����=?�3�M�v���׍���DڳU�Q�I��MZ�����۟[{]�f�<���~,���e �����A��a�J}��	�ɟ��f�r�KJV�<I���Fˆ��D�K��H����[k�_��&֘>ѷ��  �ѥ��1�BT�s��֟]�[��?��N�l�y�j�8p��Fɑ�OWޞpǰ�+T"�y��o�l�U<<oH��ac�WW��=��D<E����V�����O[���sٹ��Vw�y�?��VzjP�#�_��M����?FC�:W��A�[��%
W��m9`b��Z}�_9#�m�����"�����A�6��f5��W��ɂ� �z��N�u�$<����;d��e�|w� �!�)R�?�yrd����8���P�ԃ�m���QN	ħx�p��@����yN�uԀ"Q���,�BT��0�1K�+��(�^�"E4������V������K=����Y��@��-�������4�k�ZT�;x��K���_�Y��#�}�%)̛R1N�>�V�B=�b��Q���S���҉�����Ζ�R��˝%��tDJ�zX��R�i���vw^D�Ihs���eϝ�"�U%��Oi5�+�-��7G@$X�*��qPbA#>��N��sd���T��J�y�lW���O����
��%3�oJ,���,�>_�S Ȓ�h��������`��p��r;�|�C��E@� �z+��
<�x��~������^�D\�;g�\�PAG��pn�ژo�(����UTᅣ Z^dU��soٸ`����[�m7�$����u�����&'x]�Aϯ@ ���>�~�g.�� y��F�pY��1��۔/���W/9�xj��Qh�Y|��,�)�5Z���c�ErW�He��o�;[�Q�@0��z���L���ds�ȕ�#ϟ�߼ V �Jmt��X,:�ŏ z�+�%1�m�Kj`>���jf�A��"K�ɟ�f�k�l��L����n�v+J:�>(�m[���7�@E��D6��c�}��*���$����t���<F�Z��Żk�1�S�g.q&}���5��N/�A���ER��L5rPT����4�6��t�`��o���"�a;h�����n;{N��)A!O񁎌W/X���?��/�4���q��>w��܄J<��zFGc���f�z>�Djg�n��\��Qg�H�k�C�I�zm�h�&��m���8�heR��D�Vw���6ȴ��Q�)�+*�,���wδ�ɰ�P3�R��#�F��S>W-����=`���qc��'f@0S��_�1��7��1�bs�/����%����(\��[���_\�ҞKC��L�&+!f��h��(Ҡ��-@�_�h��U)��]�Bb�2d���c��$��`X�R}��c��"ENL���������,qw�m��^�46|B�Ni_��J����fh8���VS��u���!�K>���j���&�/��w�D��`,'~��2V���Rɯ^�_�W��ه�V�C��<	6��y�cKtFnG���{�<zvwM�r�t�[�G���P�v�<E������1x�$�s��M�<�����Pu�m���8=G�1�w���_��}�ؼN�%%�%�޴f�2i!�h�~}��i
O_px¨�9�a�Xh�	\�נ��6�1�t��{��l�\3t�x'I.t�ؙ������A�$"s��4����
�찝]�>%�,�ݣ#�4�=�,�2g���Ö?f�k'R�A�*e�~���i���+lV,��jI�����8PC�C��j�\�>"�p.�L��Y �̯{�薴Ǵ�&�Ƴ��U���
*����O�l�~)��|�Sǃ_�,�^�x �C=k{��.���5��w��*�{�8�����U��n�--���#���u��N��<�No_o����T�_R���!�����T���S��>��T���]��B�~u��D�1�{��K%�|�T;D5�Ԛq�+% �X{ISpw�7�S���Tɺ����bP 7��8Hto&�����EU3T��+�|���T�[������l��I
{�d���R�Iz|�.s �%������ja�m�N^j���Ky��x��^*+bz�w-@����c��fP�W�i��p��t�D�D|.�]�sPh����8�a˘�8^ϠЄ�u(�z^��j2%�O:��\6.�aS��q
��K�;�x化�;��a�V������ɯ�q��{�طHa�Z�����"��"r(�d���t7ݚLP� ?ч�4�j@�⋮̄��g|vীN���f�kY���h�@�D�ny�) ����J�MI����z{(�
IgF΢"�ƻ 0���S@!-PJI�
�8�,
�)(�S�2#d?#��Dz��K�p
M^e�ѧ��GNZZ1E��t6�"ts�y黭X��b�OgTu��T�T�Y0p�m�G*0
< �B�]$8w��MFIJ��;m�m��>M'z�g �s�DFƣȦ֮&�'� ��]�K@�޴��P�?2���c:���b��cѫ4L�D\æ�H��s�M��%��fy��!�1���43�"���֪�E�ZT[��K�~��������ӽ�|yɺ�)���R~_����B�7(����H��bv��,p�O��6�ɍ��z��	wp��Ş �7Շ�9[��f^*���?׽pn���W������X?DAe�d}~�ǝ��]�U�R)议@u�D�o3�P�qp�d�^��I���MIϦ��l�^X���S����.��33���>[����zFB�u��_Sgt�]Ԗ=��p���+�&y�B�� '�0U:*x�u��D���|�ΦM��}>,ȍI�-A��z��L�s�X�S�%g�n����_!���N7�m?��e�����![#�7|��oY%��1Y�*��O�w�w�P��_���~���2�1������=O�Ry{:� q49f�B��d�^v��LX�0�SOn���$��9A�;���A̋�N�+TPFLW��Vik4Wt���>��n� ��@a�R[�L����eG�8�_٥B���!DO,,�2��!C�r�f�?-,LQ�T=��Q�b�@��Ӻ�
Ez���I))��zM��ƳO�T�[��CQ����f���,\}e�%�ȍB3�lE,n�3W���;�Ej3$m�O����F��=�n���������r$/�w~.i{à@�<Э�GKu�Im�\��i+뉭�r�?�4��b������߾��MI]#���0s����c��/�7A9����[wsQ�ˇ�,�2	*m&,�֋E� g!�gG]�/����fY�r_��Z�4D�J�\��&9`����U�?itYN6(tl{'D�.'�j�n�}_�H�C��?�p�H�.c�|�S�)�P!�\䱸;dB񯷣 ���S�`�t&,´v%s��h�{!�A��h��r0т�*�`�Oc���g�	��� �	bU0���Ѭ����!��e��cC̸V���%3�w/�*�x�Q�)Mo�R�k�_��C�D�-�P���I�ʬ�諤�H.!��{���	n=����fk�>�J?Zߧ�	��	����|��VU`�hA�8tyl�N��&8f1-×QM
պ������}��w�b�}&��tq���e�h���2&��k��rV�Z��0a������7�O	��x���v�џ��=�0��A���>�14���H|)Ya4G�3<S�o3t�7< ���V:!yC���Mĕ2�����2����!����E��Ǒ3k9%V�;&ÙL���[c?Z�B��zg�g_�6�<�t��0d���|�&`�cBޞ\s9�0!���Cl�m�P~	��̀����h�,���6�@Xh���8G,\(xj5E�Y��ӄ7�P?S���	���!��mćw���t�G{B�i�g��#7�ӂu�]�_Yř$ۧ'��̳�2I��_!�^I��8��@��!	����7����Z������m�lH�OM+Af�ƫ��!s� !�<�D �ʭl�ҕ੖�b�:_����d0�d��&��|�g��?�h���~5;)����㮔��D@�u��Ӷ󷘎q֮Kj94t`�F�P	2��y�^��Ŧ�Rmw�iOp�O����S-���ڪ�]���H.���a���2�{����6H0L(�>Y́���9;׀�`�{��GG` �?���GG�j� D��.���\���<M$��
y�x���ϒ�Dlџ���X��!h0��!i��]�m��U��%XtӘ���]�7���J������K��}����h��%_��� ��?*�?$L��_I�A�4��v����W���@q��]]��K����G�"v������\��W��&)y�KP�������
�"��l�G�_+.Oa՚�U�Ϝ���?s�g������ ����r�������eMC�PK   M��W�&
�G_ �h /   images/56c78dca-afcd-4253-86bc-452069e6d2d2.png��;�_�?��h��EUKko1��Z��-�=��U�vk�-j��"�Fm����;4�W�����	ߟ�?�:��̹�Ν��8��>��~��As��			�M5=�G�>���Oz��?^7 z*$����$/Ԟ@A��ە�q>9�c�F|�Ɔ<4����ۉ�U��:Ť��ɳ���kt�4�6����Eu�>���c������P �S��c}��1wo��P޸Or��f�$�i~�	=���;�
=	��(2������WBΪ�7Jv3D�>=����2cD.����g람�oJ�{ez.��t��7!@��((��-�c�?�ks��3�?��3�?��3��߼�=R�p�������Q��N��Y���J��o�{��Z(E.kǷ����c�ٙv�kG���g���A���.}�D��Bt
�`>>U~K_�PNn����:Z�q����F��~�����{���"�'��r���;�.V�ڴ�\kM�����'3��}��wr��L�k)�,�����������������1�@��鸍�U���\�p�iY�����E��

��/���{������5N���w�0	9�U���%'��oq���0H�rrt���B=`��GCVg���
ccS�,���{o���s�����GҷNd6�B��������i4*?��:�/�z���ݹ�Ym��O�q�n����oX�loo ��Ft"�\t������^���5����R�\�&�v�Z�`WW[���Z���D�����w��˝�Zi����CO��e^²�'�Y�o ����u�`7��&_ȅ��%��%i�X�S���I�E�xMGV�*s�r�t��U�/wZߡm��Ae(C޹*H��8wʻN��>�����,G�ݫ>�!?����i���`�zDD�o��6���1�����?T�����VP�~�>m�X0��U���-���F���
,5��3QJMNQ�iу��ǽ����)��}�9RX̩�NQ�4DB�8ܗ ���2�+t!s�	
!]��3�s�����x�~���s��pB?�Յ�2�e�9q��6Fq�*����r�:;�B���.x����|>x3�_QQLJ���9w�Pzhndji�{nQD����P�f-_;�/f�H��\k}4�}�n����$�
���F~I�O3އ��<�w��OXhyzM���=Vl�\/��?;��L��wv^!��5V�F���E����T��:��O=���s�/h�cif.=k�3���8:_Z��~���r���p'^�FߧM��^�e��;;er�

㔹����������!^
�Lb���մO�{|��`����ૂ��7h�}������>�R���Jح�?ܫ1�Bo�#cTA�:<rڞV_��H����]�*����K���6߼L_����D�hcjZj�7�EJ��S�F�*���WEeZ{xx�dk�����r�6UOF9���/�%q�z����݅8}���FX���2ϗ2���j�D��:�[7g�C��p#`W0a�g$�u�U�(�߹������e�x��?��w�����E�#�S\F���d��xM�͌*��>����\�6{cc��N;������R8���/mQ6>�$ɫ@g�����k0oU��{���T�Ta�_2��(�<��Y���ogF+��!
�f��w���!� �ީ����W�kҲW�c~t~i������p�<�F����7#*>#�ϊ�_=Ŋvv��􍌍��	'��]g% .z����W�Co��zT9�O/�{�/&��7�.���H�:07E�M�EG�̔�"1	Gk�9�HI�}{�n���s�۹��Q�|t]?�{�Z~EYY~�Q�5����w��&�}����٬Us�*�M�k�,,�U^{�
�y�Ms�>��(�z:��ҰJY��<�qu!f�]3w���4'T����7'{1m]� �7t�A���jmd{�v+������]S~\`���7�ò�3F��9�|�_IJJ��$I�j��B��X(�Yo�cø��ȒS�Z1�uo>TL�}����=ˬ���nt�Qg�0�d�;La6�Yk뇋~<��lSŝ���0�Q���_Qw�{�!,���-���9�[ª<i~oь�=�s�-r���=�OTU��{�jxX��Ddd��O�6�w�4�K��<d�<��Y`�'���G�R�2����0,*5��Kf:�E"�.	��O�J������?c�m����D��\�jr�����ݭD�fF).6��en���u����ך���c�$>�E��i�ǥ����.��ψHu��tW%�KC��rZ&����Ѳ^*�<n��o-`��;}��w:4����CS~i-�4�}�B���רQH=��%%1�s�aq��^ݰFn� >���:��O�鿓� ���~2cBɸ����k��=�s��,�'���yi�\�n��~�<����>)��;w��o�>+O�:=3�nП�G������bk
u����/*G�^��`�w�!9�5)B�M٘\���dQ����p���Ⱦ۫6jQʲ9(�$�JLjD��kd�l��T�އ����gԊ��"�J��Ԃj)��E�|r��^�s

���<����֮��t6i��K��.�(�|�J������g>=H�嚘�U�t��)� ���MMM�PA�*�U��o�><�� }��w'�753�J����A�VR^>K��(z����Ut{i"Ҧ�hV�P��n�`-QIJ<Q������#M�;<��;y9��*	��FÝz��M!{�mJQ���!�� �_�'�shʋ��X�95{*�1���Q�a�V���wJ��#V�����s�%���lz�?3�o�c*�)/�|�sb���}6�_2OH\T�lQ�g����ә�2eɂЋ�A~��Q-�U��]<�A;�̻&ǰn�}M�,��Kv������ں�rLym�w֟>a�����N핂���:[@yC}Y�yMQ/��|sf���Ia�ϋ���w&��0�R�`�rמ"�꣟n8�΂����Z� g.ٹi��^k�{j������+��w�M<HC�E*J����'����^�M<���N���;�CA�ڋt�L҉[�k���3ޢ�n��L5}N-+Ē?b�(G�b,ϗt�GH%��t���?ߩ���9V8���-,��%4qu����U�*���d����M�.J�	5G�[�8yo� _� -&O�=��T����_z��w�q���g}�)��a�H�Ix	���M�jW��"Ê�k�uU� "&��%�\6a4R�)�,���¯u����+?�Lk�m��FP�0UO�al>�B����X�գ\hQ܌!5��n\��O+�B����(�i��|�7�q�����g�A�˷��%��/.1��]G������4�&������ύhP	�|��/��jmء�O>� �5XE�y=;�'߀��Ix5>��2TלTީ;G���Mxd0U��5�r+��?�`^�fATG�C���ܳ�.##�&N��}�����	ث�̪\���,�Gu��h*7ݱ�S����������I��ս�736�_o�=5�	���vE������{��]o7��G���-��ǋv��ݷ�_1��u2g��W��I3CӻnS�3\k�y�Mu�5��s2GD���/��ï���Qt �<��#�����S�'R�-x������kH�:���ژME�VNexH-H˒�Z�	1>)�X���['��O�鴉���f��q�r7~a:��y^�k�'qn-`Le�,��#
kp%~x�ѓ�u��#x�h��0��&kC�8���:P
�����J��;h��PAT�"n�	����=y<��P�ѦT��3�Garrr�W#���h{I���椦$�T���*	�~j����Hw33��,b���4�az��:7M��d�e��
���ײַr;�s�߉O�m>�h�u f�@(G�#V�k�P�xB^S4mry�onaʁkm�� [�56�.�����5d�n�5�t.��lj �rj ��]R����pHq<�C�c�@���§xSq�h��y���w�n����>O����i���Ĩ%���%[Cl���Kˬ,j���z����jvV�k%k�)IW��sާ&�lV?��z��:s��X8O�~�*�m5��6���O�vf��S!"1{?���R(J�6��G?�ܧ���C,�_�->�	���� Iw�ZM5k��-�`��q��r+���[��nQ�D�+��h�A99򂁛��D����!z���G�q�Ι�T�dөZ��v��$ �W��tj]ĕ�6���;%ͫ�ҹm��D�+��c
�t�w��
���0������ZE�E�q6+ZP�R����DO^�����������1��i�gL>����4�Rh�����\b��U�7˿�H3a��w >��X8���ޏ� y��[W/�������a�&�2��ѥd���N=������>����g��F�n�KI-�8W����Y����0��f7�����#d��!iZL|V��*F$���V��o�D�bJ�o.��)���1|`ģ��w�YH�M	M��]k�n�i�bgr�~���S��������q��t7�gE��0l@:ߺ|���@���j݆��C���g�I�5/Y��v^zJ�9�����a�Mf������_�_^^&		���އo���L:�鳃�������1
�q�ix�t�|�OR3��F��N��[�+_�Y5:���*GX�� �BqE���n���]߂ό��7m� ��=;O���l�g~54<s,�r�*^��2�tW[8��fm�JO���!΁aO�'��'A�����L��j�b���8���#����!��=P+L�^z��>ۄ��ƌ7tP�N
��O��� �"j�v::�����	Y�L����a�H�d�T�g��L�G�ג��<�q-�g�kk�̖�)R���6G	Ҵ�:w�/:����2��R�@������}�Q^�^r2?2
u~�aϹ�?�L�}�d�D��_�1b8�����2!V3!��Cq,�&W��+)��h�󰔕?����Ly��G0�\��g�����կz�B�Ҝ�o�CԖFTA��P3JӢ��*L�����|0�n�sT9��gߟ�z��GS4�I�(`a�+:�8�G�	}f]�����	beE��t�9�&%�OVX �_i�C�C�7�>�:�{��d 2u�f`��_�]���k�]g����|7��v�v�c�͝Ϟ(+��(1��OM].o�M\�۱�`<�Y����'#?��f�y�f�~fW����:�(�UT8�MwԸ�5Noy���05���{,��Y���ᬧ�i�/9�$�R<`n2�� (�t�����v�FV#��ۮGb*�+=��.e�RW��u�Rm�s�H�hB1��"
��tw����Σ}ٙnm�&�E�#4d�C޷T^7)���]8!U8�]	�J:�L��4g�qA�#��|q��T������J7��m-�66_�K����jp�|>;B��-9��j�g�Hڜg'"a�s�L�k�/)���!����Z���ApN��榫�C� W8_�����usP�U�)Ս~k��ϯ�5g�;ڨO�����_<�nb2�	�|�!�߀�<��9D�����(�;4��I�;�Jha����f	�}��ȳ艚�)��l� �9e�K6���X�0�C��G�	<�H&�	�8W| a�`˹N�R�(K��&�|(���ѳ5�壍�%Y�>kY ¼��)��+j�L޽�u�-o� �M������ҝgyo��@4��?�z�fU:|Th����("i�GW�aEΪ���(I����3L��t]2[᰽߈ӝ������?)`���f��y���Z������\��E��4� W�������vM�V�\���wð'��M�>�\�Qqr�n�_�ֈ�Ƶ
��A��$B�ěҬ��J�@=�2����y̺���2�Ó���A���f~RIb�ɞ�'�+`����J�����3��ͻ�>����g�]]yRI8 ���, ��}�:�҉,���a�N�-���Ût�0A'M�B2�ȵ��;, H���ԝoVT���O�ܹ��)�.aK�q!�>Hgv���N�\�k[�<fQ��Mm��V��Ø�C8���$���B&&[��T��wW�u��m�]��WD��W���C�DN/m�垞㔮S�kI�vRzǇb�s�(i%��a��I��>LK�g�U�`�γo7���4M�]v�P�����xJ��E�=a��N��Sh�/���?��-[k�u*Ny���q7���e!��6f�x�`BC~�D(����ԗ|�m{O�r3Yf	���&�N����L�7I�gUYf(l^)�p���(S��n*Z����H�rM�8�����{���BϲZ�[�9�'�L�V�\[�q.�$x�Zh�FU���X�w�ᜪ�i1nɣ��2����qf��S��7�xA8�<!���e��?�b�������-��h���9��\�f���hO� 8dK�?��y-�;og����~���U�K�O+ze�r��q���wU�+q�Z�5��b�Z�;éU �Y�ǻ�#��꧞�}7{���iKϮ �E�kkL�Ze��w�-��;[��'5�ea�E.��p� T�f�f�WOߟ�7�KzH�tr��9�O =������ ۵�C��C�:�bB����m�	�ƕ>⚋aő�ܨoe���ܢ�	�l����	AZ�?��\���k�8s,`J���ǵ���X��B�� ��Y��:S>h1:���E��.R��M!︯�w�(�o��K�������UY�8�M��?��n<�h��]�����*\Z^���O�a|�ʩ�GS�'\��̵��͊�2�L�cMĞ���K���x�p9���i�y�oL��y�k�8D�֤r�W�i�={����ƼdAș��UHKM�`]��!!5q�X��|���F���Ws%�X����JO��|��6B�&����~i?�߲E�T9YG&�),�r����bm���d��<̘��,���R��J���[�, �7"l����Ǩ�_R����m��a��J�cȱ�DN�"ڛ�4�@ȥќŒB̫D��5�a1tf���*7���p��c�G��l���v�<��f�d����l���*��AW�N_�)��i������x�3v�x�sI+7�vww����{�>���>���OMNu4Wg�NRn|�^ҢM�V�����ÍS�I�vA:hY�jj݂yc����^咱��jժ��d�v���K1�:�߹�Tƕ�$��ȱ��Tֶ��*;aY5S�A���(l ��)��k�S�Oa:�����0~ �o�@ �3E��Yg�@f�Y�5dh4��k���IBz�ۏ�^��U%�q�����W0��� ���e�^�;=jp@�%�*m�H R:��GYCc���y�Qr���GD��cS��gs{1�~Nߊ�sN�a�k�r���J@jMFb)"E��_CpN� !z9��6LC��C���$�E$8�Z����>,($u���?�P:~�{�Rk�sq��n]�3-��ࡲ@a��K��A�$2��++ۮדz�����_��^�q5���q)�z����"e�kIgg��u��-f�>������=��BչׯTW&�(�@�;��]��6N�ݓ�s��z/#�r�>ž{8���U a��3������K�q 1N���FF���Q�����Æ3>�-���b=�
��N=��O}H���j*���M�2r�w6S�E���A�Es=K[�~�ׇ�ټv�/�~�}fk�H��^��Vc#ځ�xp��e�{��c5]�≬9��J��p0G�a���k���wC������I��d��!s�!�^�d�A��Ϛ}EK���������!0��S�㗖ă`B�p�Fh��rP����mZ	xx�}�^�c p$<y82����&r��qg�ړ:_�\gy���
*lt��¤!���l�^�E���8C!������H�!�,��/?�%�Dp@�k�s ���^�hYK/��{%�e�x��(QK�5��2�:�$��?֖J���w׊	RtL��E�k{�9|q`��k��0���I2������H��84w����c@X����I���}!D��u"��h)`smU������XD�lg�D�L�ƥ� hs��i�vg�$�/��Z��N7]4�e�D����V�~Eu#>Ƀ��6���#��hR�WN�~%���K��&|e#����j�$��t�����o�a�q�i��;;{�u�����Ja���f+C���_�S<m�u�C�q�l�e׫4%
��>c>��f��@<��iZ>�){�����H�D�������Z���m*����s� >p�r�m4���3���lV��e�2�s��7�;ݭ��+Pm��̊S?��]+8���L�>����L����U!_035���k_��6yXፙ��5�YY�� j�n�=���!�*��e�_r2�r -����>9V�s���M����yjj�g2�B�zݬk���.�ﳧ�.��Ӎ�{�KWzA��j�0���K6m�EԴ,�M5n��y��N	
�o-���N�IaZ��������Q�3R��S�ө?�7C�T�S^h7|7*/媐ښ�A5������\��P�i�AW�-�֣��4֢��3|�c;��Q���X����
�ViZ�z`�eb�a�9�3�+���ſ�e��L�X4��3�I�c�UVAnF��wW��OF)��!3#S?��pSb��ZHH?p_�B)�i��@�1�aY؋(򠞍�� 7X�_��Г�%�j��OC�yw��TYr�n�	������Of4��J���:���N_8$p�Ų2�3n�N��Pfs;��U�l�PÁV�P�`���� ���OW�z�>�>�dL�����g�~)%ԅKʏwF:妐e̼y,E�(��tS���8Q�4�򐑿���BG�J8��머((T��/
us��(���k��c��X������/O(�&&X�Q(����K�'F�����W!ε бo��jT��Ñ��^��5̉;��%�5$���+��h_��b�h�c���!��y��'�X_���3e NOz���-Ae�+Ḉ�аv��H!�-"(.�X��6r�����3��h�,&nۀޥ��,�
�:��|���I� cQ��ƌA����B�b�,���=1k�=/ള/t߈�Ip/�l�xZ�}�Q���m�c�=��s��1?�_ig�mU��짇�8����:V�o6�N�3�8Oj�������ܟ��-�kq�8DN�����p��'2�<���տ)��9�_"�����h���xC��t�x4W#��F�w���$͵��8�:b�?e��{�v�=�w�iY�I�����c�mK�~�q���K4��m�gu���b�W��i�Li�ly?L������,�Υ��T�4�W�l���精���z�=����r�.��MV}x���Ӛ�Cȁ^$"2zMn��?�}���}�$Dk�1�x���G!)m
�Rڨ?@�(���T�[�oV���^�Q�8M֮/�Mm��G�"^��i�]%;�8n�,kC����A�ˁ�FJ��c�r����L�}����H����z���!B��;غ$�nȝXGdg����jH��W �z��
�92<Jm��v��`�]bq�ώ�d�`�K6���ͥ�X$PvDlHޙ���f�}�83#C���ڽZSM �Y�*@����'�rT���T�WtA�<$Mwnư=��Q\}n��YZm�۩��i4�Y��KټE�@��_�=��(��*��s{v͎�BӞ�⣋S��K �-�ך�;���u��M�دڷ��g�,�P��]UB�}X�z{�*�R�.7\�[���o��wpǶ��4ߢrS���4[Q��Rr�'�����{l�cŶ���.�Tq=�k��YS2�K����x��C��4&M�x�#�f_�� &�>��v�j��My�����MoU��}?���7R���a��gX�B��8���,��i�3VN5~UI���d�6������YgqB��O��s�KDe%�����7�17��������������d��)T�1<�<��o:H�8��.��M��9�L"�"�+�a��.va��1�S���Ư��@Q��b؝8����ݹ�u������Ix:�'�����x��s�'��<�Fw�,r�ZM�5�p)ڝ�/�x�z���U�#�K{�^K��Ѫ�@,QViNg�ч����58��)�>r���r5K����a����"��H�J�Eϲ�Y?��ر���fjAx�U/�=\�I�a=�$qNi�E۰Q2)��;T�g��&i=؄��e1Zr�КoLf�/]�4ȶ�M�VvES�6�槦�3������=CsT�|��v��@�/������@-!��\�yS\�,����r�#�A{��3����!��߷1<:�dX����2^_�S��ٚs�a]K+rkMIJ!2����|�o�|.���qMDS3��O�oy7������[V�% ��������~��\p���jQ��2�����Z�C��mV���p����E{�;n�?Ƀ&���a��gXyy�
�I�>x�4ɵ8	=�u�Z����hX��� �4Jz�M~4��ɫ����U�ր�T��υ{w.ڤ�-��j]Aq���Ic���:a�~ng!�Ug-f؋+N�<�*�2�(J�������UF�}�4sgW]6�"T-+��.ϲ��f;`&d�{/LG�2��K,��S�0�a�O�GbGA<ʑ��ɵ2�ta�e��5�����gk(�	�<8[��0����~"FV������]�ne��#UiWG�AQ�/v1��@@�d�DT�^��#˅*���v\333n0X=��!!�W M}�XC�����V�* 
�`��Z���4R�m�!��=��~��5��G�V��nf� �2ӯ;K�<&��_>��_kN�p<�W��g����O�̙��IР�q��������_���!�b��L{��ߙ>���+�Ñ5Rw��P��x��ޡ��0��ʈ��)��*|�[=�7#U51���R�Uh�NК�������J�*Gm�L�u��J��޼�xsǸbځۚZ���V?���ں�ß���N��9����r��� ��-I�&A�'���Rm��י���${��W��t��n\�wgx�������h�l���\���?���7���m���ui{�Q>��Q�si����AK����_p�e3���G�Z0]	�'��������i��+(�d�����H����J��F���G��ְ@?,�e�xu�'Հ L�}�=���mf٧�7l+NX������K̽<c�r`�˄�8��Bn��'��|9��m��j����?���Hx�*��C��1�y��������)�^��M2*�v��|�o�7���?��z�V��,�I�Ll[_QRa�?�l�4�9�!��Ѕ�u��B�
��F
�e��rv2�OJ�Y������w4�3��>�353�L�j?�"ٳk��Nt�+|���iYH��i����ӵ^OV{�9��/+2#��øv>S^H'��ą]��pSN��xP?�D܋�z=N�MhX�p����B̦7~����`�+U��6f��n�������RO�`J_eL�`�؂d�{��ߞX��3.<�߿�ŗ����K�qY�.�i9.-=?�*���3�(�0-L�?4l�=롺�T�>�����$��eߢ(��,ʘ��۹�vQ�rk�Hѕd3+&��u7�^��ȭO/�Lq����S��g�s��]xV�U�m�]�!}�C��%�HhF���A���96[����8� 6Io!�^�_��s)ßE�Z/�PL��N���Q(��-8�ޏ��Zj���ʉO�chI�@`��
���*��Y�w&��#5�|��#"�U����pP}P����(��CV�tX`T�,������nVw�����'�94eqK�5Dz������h���2�l�p+��~A7��^�e\j<��V.|�N!�`��@����q�ܺ��� �&� �L
H){�(-M�WH@��9
g�x/�G�F�͐�G�d�wvv������ъ�e����7Z5{?�ƥܒl��s�FFb��T͚n�
O/v�&\���|�C�&�Sq�qt��`#� �Lt�� �zǢ��3�����$KA�}�ro�Ψ�5^�w�G6��-�g�.Ǐ�ng������K;��
�q�@��(���K ����,�ѓ#��z��'Fu)��F��霘d;<�#+{����$Fo�滠�y�gY��䆒ɢNiR��ޞ��u���,M@�Q��Z���f��,oL#�L��ӭ�����.86�m�O ֚�?�m�&��U�����}/������ceɳ��SMx:l���,ql9a��e<z��q��c����@]@C�-���G�)ט��'fRkͰ�����#:�7���2��2�\�c�Ӝ������Ƞ������&�uHd����|�p
���%��aɬz�$��M`/�&K�AB�z�|�'�4T�T�t���&�?��n���]�:�Ә��z?� ���]�'�UW�vUN�6�I�Ё\ʲ�����D"�J�����bvn�����N����}�˷�zc�V�Kv���� 1O
�m����I r����-�6��u?p˷��*6�W�t�<��u���uC�����D�⌫{��}'h.�I���rҗƆ:�2V.װ�*A��n���x��c;�7j�/ ��V_hxn�l�;!��N ���$�2��AϥE$ �*�p9�
:�H)��z>=��U�h�>�%Jo5�/?m!�����w�%4ۚ�/ȼ~��O�R������v��R�~��Cо�sqpWL�����7�6,Wt0Q�&�yCu���:���M����,c����& ٦z�۟{�h���tnUxFܛ��@�ۡ����������V*�*5}��Z���Q�)��p��%���f4ޡU<�*E�!!׭rg�u#��+��z��8����>�Z���tm5�y)hp�j��ۯ�=��5��4>V�Q8x��O!�L�S�N)� ��8��swu<��疉��x����}'��يMk=\x�-|�;��jR�b�6&����qM�1笋dɸ`����f�d����o��V��������)����,��N��Z�觇olo|MIj�����������C�έ��h	*��V����pQ\U��a�QJN,���Tejj��2!r͡kۧ���{����3�ξNJ�ȍ�>�P1w��}����J�
!����)�-$��M�����ڡ��1\�;�5>n�M.���Ap81�b�e�d�~jb�E�ߐp�I��O�]�"B���u'�V��4$��|�����N�G��7Qu{�-��"��L;�c�� 3��2Jh�jT"b	=�
�?��~�K��Q�5�j�+���yÚ���']rl����J�Ni��_9�����l_���R�eU/�O*�;H�u�\����AxL;��v��bEl���T?�DP�>7
p���m-��)5���+A;cPq&�M�>��L-BӖb[�:�c��n���k#%7ů�/����v4�ިf�!��	qm�c����8x垜�`c퉡�,[�P<��5-Di `�s�6���}{r?��]J�Z��(�����]	7A1{K�,��4i����$��)R�d�ޓr�[Ԯ���ц�Ԗ�K�R|�����sU���&�-(��C���.��?I7C���o_T�4l�7]�@2�Y���cy�:o/Y�����Zmh�O��5i���Y�@��u�jZ�	�nyZ� ���'��{S&a��s��1�c��R<=��#�M^�^��3�%U�u�c�s+�d}W�r��>�i��ffb�8�`��c�1�s⤄W54z�e�>l��i�Ђ�D�d�!no���N�0Yg�˧媛�ϱ�Lܞ��6���=^�L���ጂ������c�8�5�����i�ݿ���e՛`P�,]f����H��t�܌BT�������N<�_�^NP�'~f,����P�*�dl�����D�@�`g���2�h���o�L�BC�'��{u�+��F��˜���O�]<��9>�Z�Jco��w�%�:\p�0�3�B��Q�Q��d�ۄE3�p1 ޥE����ߐ }���3�D������_�Ou��m��޴!M|G%F��o�D�"�������Rx��IT�)�ۆgY� ύCഎГSG!&��Pnj�=/UʟG^	W$y�}��(��3BxRY��>�����A�yA*�-"{��9D�^��#�O��U��C�FOihߖF p��̉��]��g+�����h��ɯ��8�y'e����ճ��B�|���ܽ7�C����Xi7�n�ڮ
�\��zY���ɓ�l�:�����B��:F$i�E̚�PB��.�g�@m�C����-*/_d�[��ֹ�X�N*g��
���9@��O���������~�N�M��p���N�C�F�g8]hV�&���~��-�*Կ_ �e�d�?�)���͗�_�;��<���ma���@[lR��E_��B��F\|��w����[l>7++{�8��.a�U:% `���SO�<�_S纼����+�]P�ʠp��Μ�������}w�P7ϙ<���L�LvΕ8&�8c��IšLȈ�j��j�Bj�_�d��?�5s��h+,�u0��l�#l�)�Ҡ�,2y��=F$�z�i"��;�$T����6�5~�u�h=����-� 3�E��>��]�f�����}ek(�c�����p��r]�����A�p��_�kY�MR>qM���]�_���j>󝕝w�|����_��u:��f�(�O<�V�^���pO��t��m���|�K���T�f���1�C���H(!�ט�]�8UF���1�x����-Rr����_-�A�� ���=<�Bw�p��ox]4�ck��"���J�R����fō�K�\�\��+:=������.P�s'�C���>"�9�֏Ե33ɏ��o��C(� s@�o�2sR�=pvu}�6B����MM!|Γ���:O����D�.��S�G�"w�,��o������K��>��J՟�"f �6����ooHp�{Xx�:�3iϻ�<vf��dVP��E�|טL2ȁ���} @��!Bs�~_+ɴ#S[�����K��WWv���'���p;�����C�>��fƕ��O�k��O#�~���ڼiҷ���d�`#\�oFܽs6"�y�΁������?Ce<v"��/����y����z�<壣��ϫ�� �^ۧ!��7��*�a���FJC��kG�~���)�C��:O�s�P�ȟ �������Cl���}�^`�p�[��il���C��W�'ݹW�����f�*��g%��YiX���9��1Y��Z���R^�����zW��.�Z��2��{��&��K$6�Uj��&rr������qs�����hR����'���������5)���ۭ/Zwc4ֆw��g�\��	��f=K���Ĥ��L3tYXۧ���������ӂK/�sw�-L�j� �w�$��PS����jw�l:u&Z���@v��r��l�aL���|�1R�=%��O�3"�Yr��:��s{t��1�j+�������ek����h6����gåU`���j	�����0�*�*��'i��$��-�𱭥�L��^�\]�������F?�*�`a���9٭��:*0#��]�gU�>���g��(�t=�S{dTGF�U��� ����Ķ^J}ӆ�m��w��_v�n��%��˔��k�d�)_��h;<���S��u�oZ^�4��|LAb5�<����*��+S�O�",_ƾ�z��Ϫ*{ـ� '���������6�zuA��/���8Vv#-Nvq�H���4&���n�76e�e��g\�D�=b�Q��V��i��/;�gQ�5�Q������o�n����O&�p|~���PEF��K�o���ee����y���J���@�'�
grx�ţ~յ�Ɇ6�	�ւ�ݴ���{�}��O����2��C?]�/�A�s�M��#^pJ�~�s�s�;
52�T�6��'�&�,2�'�1�}��&_����pv�١'\�E�&V���,�s��3"��~yF���z-��5�]D����M0�M��̬��W���&\/S�����Xyn�I+F����9�	F� F@��׵{X��FF=gMą�X3���t��wZ(�� u��ĴE+�I��D��㣯`lԍk�R#��Q+������v.6���ӑc'�@��]DV)��Υ��_����瞵2���������BBL�P�ۧ���)����fD�>L+��Na>gN���8GD�yA���]ק�z"3|h�:�j��l'�yD}�F'�� ��FQ9����ȶw����^�k�;"?�Q���P� ��>����Ǟ�O�����-eq�@ xK���3KW.�W�k����?ƮR[�;�VΑo���ސ��O�r�,��-/��c�'C(�![�Y�Ʉ�y}a~�LAFu\�]rQ�B�"u[s���%*OT �s�6r<s�f#\���^Qae�³
�R�̓�˓�ܚ;8���1T�R���G�!Ϋu �$0c��l�&!̟Hy�v���r.S�Ĥк�	�+� ŵH��';�mlz�s6K��69�׏��� h�8ڃCLۗJ/����5O�N`���	Q�:���Gy���L<9d����1��l���2�2�CԗOO~����}&�����K�G�v�T��y�^�\���/X4�._��.�[n������0*�C�����5#[��0�Vm^�_Ǐ���
�u}��!�ԇ<r		��`��
�c�a|���3��%{�?2d9��C�q������#��={�s��?074�_��r��+���h~lgggxscە�l�xв�Dati���]�c%u��Y<]`vhޭ�;�@d}�r�֔%����{�5��/GarkzP�6m�r>.Lo#���[�r)�!�˗����&�1�4��pyn�P����9k��k���p�5�#52c��{Z`��� R�+�
yax��%dϼ,�OS�C���T�i,c`�m�{gʡ������k���ַ�e]Ϙ�;J9���u?��i�"O��ᝂ%׃�j�x���=��Kލ��8טp�w��ֳ�G}X+����ͮ�k��^u !�A5U�vS�^M;�[�ӿ�)S�c���{���@e��NC���p�����:�F�.};��e�h鍘�icT���7���Li���à�;x��y	��m� �]���^P�|�Dr];��,��I��BٽO�7}�0��[�"�x����G���uۉW���X ��З�6���W�7hww7������F��B?�9�H�n�j����Hݫ�/Z>eq¼�[��M�qB��i�Oy�x�x=,�"6�W{�"2�`1�-o���m��{�/��`���|���Y#Db2�89'Ǣ�\T~x��}�H�7�k��3�){^Z�O^g~����6�T���8�����#�u
�*�o�@K�,]��b����<T��~���MfD�FV�޴�����Dk����w�ݩ�O��!�#Mwشfm}=U*��!$d�lt��������Gh��o��R�zn���޶��us��q�
�r�0���}�v��8<�`��4C�������\�͵u3&��NQ��'��q��]����l�C�_�����\���M?��?kǼ��������鬒���߫@qo�DF���]�C�[�ꞗa@�d�F��|9���p}�{��n;s��]�����Û��\�ek{oa|lxa�س����yt�O?������o�X�yp��+��'��8>6yn~a~��r{�w��
i��r[�N����
��;7w��w�9����97������Z��W�7����J��:����/n��˷�5�7��_YL����.d�1Up�ˮD>c#,��n)u�*w��%�����Y�����8���ܹ>S�f^����z2���cD9o�)�E��@�%�VW2�z�[�U�.o��n�)�����E�n"�	Ϲ� 2	�׊����=��E
(��>"�^�=-@�XQ��9���y��A�ҷ�@��5������]�v�n��&;�j�Qy�,��8V�.4����2�C��+�f��w����KܶL��;�������/_HՃ������A
���c_O�.\0�����ͭ4>9ajt���s�����_� ���M�Nx_��ǽ~�N��O=�دwK���V?zu;i�S�Ͼ�̟>�<z�;��{���F�t�����z� �����B�e�a`1~��5���m_�z��Z�N�c!|W0����_�U[�g���O��1���%��^ظ�����'ƿ��������y����_��g����r��[n���ӓ_|���_��>��6@��!��t�?��X���[G66�m!�5|A��q�a5���c�xD��2u���B�z���ɓ@�"��`yU��:�I�����	��Y(ln���G���(j��̋�6�|�Gm2j�G;��K���B��< w�"a�e������{ÞZ��B���++��'�Ԯf�I,u����eλ��3�)������fQ�������_��wN���H^�B��^��dk��5�ݽ
��F *�#]�et�5{�����������][��%ԣ�Peȫ!P�>}��\��
%y�3}�g������*�rz�{ߛ��=ώRݺ�U�,�@����&��n����t�rz��glG��Hss&���q�����{M������P��=�H�a�=a�-_�q�·�6;5�u��+ݾk:�a���@���?2N��:,f�>CڋqKx�t��J���/��a\0n��\_tmY��:�g�+��y��| t�j{ =�n�ۛY���9����������G������䅗_������'�z®����Zʥ�n9{�O��?�#_y��1�>E�M'���ݹ����~��ʏnnm٢�|kw��w����<<�̯u��y�)�\ �^1���k�iH�e�EB]�X�\@�-Q�e4d�E��;�Xƨ��(}A�pc�l�1�9)�!B���nyg5�25Dzx���8$%o��X-t��z�,U�nьL$ŢH���*�f�y���+��YJ!�B](y(�����r����`��-�MhO�q����|���w��Y��+l�R���K$�����x���aGG�y�w~n���	�,5Qt"nz���yÖ��9㽢>�$�ſ�_�Dh{��wޓy�ٶ�m�g���s'�r�\���ݝm�7}w{3���sv}����0�F%���{z^g�TA��ALf��K���~̣~�}��.~�4Ҏ��m~eD��;96n�=��K�4r���6(���E�佳���\ky����{�^���^	��`���Jv��;w��?�י/sW�d�\[��r���#�G_��Q����P>�?u��;�(|�k_9�^D�,ZU.�Q???�+��_�K�^����`Zo*���t�׮������M[�[ikw�%"�����Nl����TX�p���;��[����In^�A�|��n[�Y �i�hYP�%X��l#H��V�g��E�}B)���<�u�H�n6�ϴ�	BX:����A�5k��|>�eAc��_e{���'��d�ysi���W�K����vV�q�l��!�--�S���)!SBϊ�0'<.ڱ�q��XP~�a�2`����6CF�����;�����Cۢ��U�h�ܵ�c$�ԅ9C䜏92�����ۭ��K77�@�Dl��~���Ϟ��~��Vb�8��S�N>���B�����f���ͤC�`;��ҋ6��#�\a�w�+��0�����],�������9;~Mi��jY�wRfg�Y�"J2�
��,���_oz^��ͳ��5��*���Ra:��%U�"�7E}�������XF�F�>� }E�T�"�qro���	��.x���G-��񈂼��w��+��@��+�?z�?�p����׏S|S}}�3��q�o_]Z��˫�]�9���y���HV�a����MTfdF轡v]0���JB��E�¥�6�"'�����)<������Xhx����P;s�3���R0+��y9mEe4�.�WK��91&�����z�E�c��js��*�z���~�0.��eD���W�3���YY�8tn�&��'��g���-��c����ꊍѼ�|�r�������q�j�#��{��._��m��|Y�հ�{	��y�M#����a44�Fp���O'N�2B�د�M�<�tz�_�����k�L/}���y� )!v=3#�E9b�V��l�V�=�?2�T�\�谕{�za.\�+����qrn0�N~�ք����ȈaH��?��x��ٙ��[�
�i�uݤ-�%�*D���ݷ��0��v�i) Ke�T�]M�^� ��mL���}���\xf�1w��+2��طΈ�~�n��RT
������=�h�f�Z^��W���ؾc�(0�^������`��^��D-R�T)7��|�T*䋃ۥR�9X(���V*�򣣣����z.����C?2F��F�'�卽��^��/WVW��ۯ���k�������T6�&Iȫ��m1#�,��j�Q����E2k��yd��[aZΧNs�mf@0��~�s+cjy��ń�BJp^m��p�r�ZT-4)aX&N��$"�=�{l��w^�&��o����Ps�3#��¦<�r�:��̮��_9o�ɀR�^�����|(�zU����\N{�;����|�>�X�Q��M�����R�_��Jَs�>O��
���2����h�R�\�b�Ő �.��ױ�'��o~P��1]�v%}��0�9���w�B���f�ښb(-��_^��ZuRu�q|���/��O<�N�|/^(Dl�'i��{ь��!8#l0?�X���9�sKQ�����V��qR�� ˡr�����t���y�Yc�"65]f4�3���/fF�WJ�K��<dj�eK�Z��Pe0z��/=�h�3�)E����'�p-{ׄ��o�ާ��|Gypl���'�w+(�&�8�瘌gfj��wm��u��|�N�f�f}��W���J�b�X,�J��@�\��+�r�R/��{�����������K�c��FF�j��#�S��*C[��`ur�T������r�]ynh҈�ݸ���~ue�}W._�����#,&;����E�Ɨ���Yi�ʘ^�q�[���=Z�[>hp����Ɓ��<�/cA�<���C�,l��>�z��-��F�����yr��W�W����p.�{	�[����q06�Y�{�`�H�p��{�,R��7�>�"ƹY,y���B���cA�Q��=�0lo�7Dka� >>����|Z���v�3c�h��A�|�k3~i�W8_^�v<Cm���ڵ����M+�#j��g>c��6�',�k�	�3'T�\T�`EɚU�X��R�7��	���o׭��Z�9���5��ǽa�U `>4<���r6�:�M��-���U���7ƪ��1����À��ЈGg��~go�� %�1I����ꔚ�p�7�aj��a�Qăk���%��C�-��-�JF���<��:6⡻!�߹_��g�c{�����qq�q�6���SO�y�X���"�߷�����@H�E�R��O?ލ�q�_",��^Z��+����Yä^�W���[��y�;OևGF�+�ݑ�����������''&����R�<=>uqd��q�̙��z��W��;�( ��6����/��K�+#x�x���i��+_��5qN�Jj(�@�?��!�)K��M:T�3��5�[H���ޯqH���c๮ʷ�o# _|��X�X�}��@��y����MHڦ���P��o�E6|l�B���5"�c�,�xN�D�{�{�Y�wi�\�ż�B�L��s	_�.zC�2�X���F)2�dl@�jr�Bʢ���`:>b���n����X����{������ܳ��ܽѭ��S?�Sv�ȑ�#1Ҥ�/�À�p��.v��b���di���SOx5��T:}��ip�7�Nۻ[���;U���.�f�F��o���x�w���T(�-�O��ݸ��Z���r#��u���N�ci�B�e�R7��--T�۵'���14���GF���G�{����)��V�;��9��_"@��rO�q�(,�24��Ѝ'v7�✟��������'����\�(J���Qm�sJ���c�ŰR�V˴�j�Qq���Y��aK�B��qwd�Hװ�� ��(�0?���P�u)�%=^�\J]i��Z��|�e �� ��@�2������������������&&&��p��S��RZ!��d7�y���KW�¥�����ni��v�|����j�ѵ�.�UY�8��O*-���\��e�vj}3B���Q�o��u��W gQ֑K!e}q�7���,F��z����]k.�g�_R9����/~�6HQ�3�cq�0���ג+�)�Ղ"4�$dt��%��~����g [س��U��������cx��TB��m+cB��H��,�(�H���AX�w��|�pi    IDAT�+�y/�ٰi�a&��0D�����	 ����o�j��k5�YF@�}��B�X6���2��z�<E�Yif¸��?�LX�a��?�þ�N�`���&�pigg�T��v��Ŵ��bdJ
ffz�{�����Q}�x��mS�◩�m{ٔ�mW�*�.�0��x̻�<t<�^�J͆ V��	�J�w�GY�M|0N�����M�P����?������b�6>�\�M��ӿN�J��s�\��p�9�PY��i��a����7-/����~D:8��>�9�_ m�5�ccp?p���[ؿ\��6�k������:٭S�'��O�%R��R߈��qO���U������K�f����:�����^�EԽQ-��g�&��Ԛ��O?Zz� \GU����K��3W'g��������#/���|vqq�Ʀ��k���N�++�;��|�jyg������廢�!�hy�6eB����n�:�hq����D(��k"��\�K=/r�o�H��_4�lE`*_��b��@<D�X ]�0q?y��Rs	��1~y��7asc��Ѩ�!q�}:)hN�M�i�˖����0�«���7��B�·�}�����*�
�^;�����V��IK�o�\kQ�!MDqDl�(;L�c�[���Sچ��E��yh�`,]�q��1ǣ��C�r,T��?�-��>�n��v3&��'�E��P(ts�l�b�˥�!߬ei���/�"����̜w{+�&+�����?���(��﯏�
.DQ L�y��y�CX�-W!���/w;�O��عg���(MY�a����V��T
�o�+�J7yd�h�q����2�����L�������*TjN�n{��hϩ������4�1�ؤ����<��L��Cx؄Ιse�Zum�9Ȟ4��~� �Q޻Fp/p���A�H�	���!2@��kF�!r�둽W8�an ��aT,ڸO"����+zc�^�Bc�}!!"���a�Y=~��G��V�7:�4::viqq�s3_>vl��/9r��x�%�+����y������zbm�]���ݻ��Yw��t�0(D{���mU���31V���/�y��eݓ#7��B�"/)�{-m����T@O����Dl��T~#A絜��NWQn�|d�[��<XT�@>�N�����}KW�^o^�V[�{��0��	���D�������\m�ӭ�9��a1���T8Y�8�)�wz��U+�b.�>>��TJ�g������5���_��<�XJ�Eg6ۖ��yg=�[isk=��/�B�P)���ݳ�pw��O	������w6������� 7R&_^ȗ��%��� &
y�o�O�iY<f!�
BA���y��"�����Ę��֖7�����n�x�ã#	��k,�F��qS~�� iR;.p���{�2di p%U�f+��:�N*�
��67]���7�q�5�=Bf�-�l�W�;i�3��yBW����)����:���1j\ ���V�x�A�^��@���s�=��`8��Lu�e�Q�##SA�x@����;'U��D��������w]�:$�UƴGp��2*\�)��â5�ϊ�e��W#,9%������އa�966vejr������;y����_���#k}�lo�I�n����.?��/]z/����-�*M��+;6e5׽_�W�93Q��VV�n\�{_׵�O֮{7^���r��{=t}	���>-",4�R�u�̼f��O��K��]޷y���+n�ֲ�Ӷ�*t΂��0��i��8<|/B��C&��wӂ���9�����=woϵ��խ����
*?�Z��ʕ����rcf{w'�ol���Q3�[/u�g§���sϦ���i~q�Ț���j�7��C1O����ҳ�\+�W!�y���f<����׫�yo�r~ 0˶���sg��{!
� �܀-�2��"�#n���@ &��Oϙ7��*x�^0�f|ܼLH���~�Y����C�iD��Ot�+U��^�2�R�+�T��>���4T����(��ƇY}z"�с�?d��^�o��C����F����N{Y*���7D�
ȣ�s�������9�	�� ��)��n��P�A�3��ܗJð֠��u��������>��/z*Mc�T{)�}S!�,��KeW��C ZǸ��f����a�F�^�Ǐ�#Z�<*�xE�j�QT�H���0E����
\���W�..<1;;�s�3�_���;^�I��6%ķ��_7B�ι��⅋;V�z�Ε/�	pZnwC��]��D��^�Y��%Hp���������Z̽!����w��@���+˹����T�-c�˦/�B�2L������G�J��ϳ0��UY�]��cR9�@�[��ޞ��Hs�Ň>==۩*d�Ń�B@`���	�,$�QaL3>�R(�ga�lq��d���3�-�`e�Ò&� ��Կ��%���x�a������:����چ����gIJ�٬Y�Nt��nvx���	+�oy�Î/����k"�?��ʮ�:�<�sr! �D$� H�9�`�,JE�����ݫ�^������^�LkԲ�ز%��(J�L%Ӗ(�9� D��P9��*�W5��}�Wմ�H$�T��s�����N �	��DO��J���2Ogk�-n�.e�t��v�eͰ�je�������� �j���;�5a|R:���������
;�����ZY$wQ�� rx_����1L�8%����t��]��@�����=?�)��hx��S��b��>�{���[_�Վ��E�߬[���y	X�� tbD���A.��:K�e��7V:��q�bT\���'%]�%Fg��۽}Ml?�&��DL	1@c����cF�r%)�|��,%� ����
`
p�PF�g>��(���P\Vl�'5Q��5���,���y*XP凜{&��K��r��iӧO�;k���kg��qUY���@�w��-�~�d�5{�x���=����6WW����4��ݧG�ImD�^<�LG�b�/JR��yc�_���[t������K!A��k���Vd*�K8+�LZ;s�o
Sn,���oZ�K
t~'�S׮�Kkύ=R�I@���:�8ו"�����ɌGY�6��cS��S���uP57�4
M��7�"�Mᇤ�Ym��II��;ƀ(���=��so��v�}貢��(YJS��::[-�������G�
�y�a��Bm�;�b0F��Z�p��z�b��8PS�@`(c~YR��бh�r-�)�N�Z&��=��2���F�(2�c1��l�)�������2kkeo�_()�x˝����Wp& ZY�Ah(���ت��~�1��u�� 1:�mܸ>����������Y:�g>�Y�Ԇ����s��r羰+R0�WY�3*��u���y��97�����xd�R T��"�#��|K��j�R��XK)��zsLN�꧱�kR	e-�^A�5��G�U����=V��W��I�p�����ew��ap|�o��+d%�������2oJ�q�¯���W16��(��ޙ�e������9�_�9m�W�ή}t����<h{o��-�����]{���w߁�l���N ��"���Y���4s�x�h_�ڭ�X@��,+v,U���hȱ���/p�#l���G`�X���X���	�(p��%�Q~`Y��kT+@K~h�a:L�U�N�E�z.�$�d/�R�`�\�[��32�kȁ]���	P�������^�}��C�`����L��ǪV���̃��qM����'?
/������Xi��;纟������)�Bl�b6;``���3k��u�&M�f`�s(�(7KL�פ,�)~�װ���{��(#E^�WnX��H��c��ys���l���ߍ�$����b$b�����|����m�ğ��� jx����c�;:}�S��o��]�)�
�x������ ̛w^�O��?�W^����/ tw�Z�t�WnS�v�ܕ:wi��a��
���'?4��5�
��3 ���{�)�|��)G�]�0w~����1��zh��r�(���{��G{F�<��	�X�Ar%)�2Aߛr�H�TL
k��ʄ�����z�Z���q<���OJ5�(_ ��w�=\Enʔ)��wޣK.X�W_�h�{&�9�~��ر��������z�4�j-�I&���֨�9G}D`��Yy���?	
�jRK�1����}!���J2�dYKpH��n�O]ԴpD��*j!J=�
�����k�w�k�E�_-	��qK@h]�u�z�Y���cIO����Zk�f��9��\�WGGW��8���߰�o�8�s{W��p����3�-�jJ��=��_7pX��2��9����<�~� K�U�5��8�;@�ig�Cq�m��QSJ��E��{�]# ]EV�#D�ā�B*���ü��2V���3�ʚ�jn�E�R�x\����MPP�-��`�/�ʇg`5�c�>���ˊ߰�b�c�����}��t_K[�?�����[^2��������{)��_��݇q������� @�8��/-.�qaI� �^m[M�g����e,H�}�+HR{�c���̩f�T��*%�=��c�Ͼc-ECۻ�y�<+������U6VP#�����N�F�N�����Qr$�Q�!W�i�uA���, �!y��mݙ��߱���t��7��+d�a���9���l�N���?��-^���kV,��΁���H�R@���`���j�N�����r���Rg��h%@��4�=��z��y9E1+�J/���.`�曼n��h'_F)�<Z`B~Li�z���$���4��y2�&)y�8�J�ѵ��>zium��t�EOZ���M�:�P�Y�3i|�s,a�˹B��pt���Ss���	��|�~J�{s������ Qw�GȫO����SX����1���G�5&Z�閖�0aB����u :�����z�{�������k�S�,��><��;�[SҢ�^ی��C�S�N_�o����	 P�; �Հ���B|�� X)�ؤG�g�z���^9�Xf�<  ���s_�)ZU����K��˪��r�=�=����Lĥ��R֕�Dʧ���ax�����e���ٳ#�B�ڲ�rW =��`3+[\f��7�����6�ߔ�D9`bP� g���� �Z���-��y�?�N���.7c᚜SQ���ep֬YGV�Y�ߊK�B^��@ɟE���E�L�jx8[���f��C��陡̄��Hyvx�03�)�d2e��ly&�-�f�������4�<ɩ���(�%y�w<y�\8r����
��X�q����e��
��h��vW�S���#<?ֆg�8y��켹s���e�b�q`?�����?����� m�0�]��5^�m&��⻖�?����dS�Jg���-�|����KZ�Zcmb^Y�
j�gY�z�u���+�=I5s��y�����yQ�X�j[�V��%��k�Е�!�_ �1�iH��V4��qR@�V�.F�c�r��k ۸�*W��������b<7	X�;��/=�?A������-�H�N֐�R������s�>ݝ�ƶ ��~�D��5kքI���|?O����x�)Β	ik�Ӈ��3���D�s
�b�GA���ө�'��	t�4?/���F�ϊ��{2�l���-�r�{�a��A�/����;��W|�؋���fX/օ�>��G�MUB��jȷ�{!�"%W����Z���F����?����GÏ��0y�T�>�-u�� ������~����#��E�����r)w��v/	[]]�[��3.�J
v�];���w�0x�~{��mi�5����|�j��<^��G>X�Z��%j&T[Zcy��磟�k�ǈ��?���o���g~]=�ul�J���E��]Ž�Å�lOI��`�pe:=8)5��1�?8#՟��J�����f2������t:]��d*$�d��s��('Y�/�w�7�@��`����1t1=�dk��S\^���(�#+$�x��=��K�f��^���ϭ�d��fϞ������o�
�e����[{�Б�nmkmm�)���@d�f|&-�$=��N�#�d��A%+�W��XZ]BL_�w���Qhɤ���yi� �KZ��k�yb��YTd�P�u$뚗U�d��zZQf�9�$��'kY�^n��b9L�/?+7���R`ܜRt��5�T��j�ef�p^h��??��v,s\�N%6«�9�)+�{c���zl�<���򾉺��~k��a+ǉ�LAj{��z�Xi&��b���*���C��  {�P���q|��Ef��]�@,����;r���sX���=c��Kl���&ؼ���<{�hLM��h�[���m�����`u�S̔`E\��M��Ϲ��=��=�OQ�b�NS�-���)
X�7�tc���>��><��� <��Sa͚�BCc�1L]�$|����~𘍕�F&���+�3»κ�"��aLP�r˰������O�2$�b�Lk�s�N3{��w��y�̙B(��������Q�9�����L=��S'�/�we����/|�/�{�쯾���K2�Lekk_E_M*�9��/=;�N/���>o``pn:��488;0!��V+�e(�q&�O0UR�������D���oh�,s�$HC�����K�����(f�Y���(��J�>m��+�_���W�~�7�v��<}�2@?x���O�<��Ç���!��)��V�Qױ�hl	Ѥo�@�_��`���(��|�ɱ`.�\t��ä���*�#	���A���DI�#�Vz�� �"j͔�D0��͋Z$��OR�c����s�5���mAm1��q5�?`�kA���iS��X��7�9���H�"��y��MyY���Z#��.h��	��ҷ��|g�L��u����ojh�ySH��J$'0��>�����l*;��5eP���3�0$�?d��%p���9�_ꠓ'͹r�����#���U�v+C[]�VQ.z�����=cݺ�y��
�Y;����Kl|�k68� �������^\���U}�uв�x��[�=P�x�衇BwO��_���k��޻wx�g,Mm鲋����߆U�V��|���O=��)D�ZP�5C�=~�Δ>Wؤ���h
y��=��D�C�w��������,3��-��򠪌^=�"��
q�#k[p��7�s>=�s����iˊ��뮻��� �m۶�����t:=���{a:�^��ݳ6ݗ��?�?m```��8�މ��9�����B	���N�|x	�w˨��1W�0��)��9��Q�.L�4�>	�b��?Y�p��su��zK }dd���m�����|��ރ���^F|�/	���^�Ĳ�E%�Z5�)V:#�I�@]�,xS�2�I�] /W�E�%�����ŋ�R~��=p@Pb$�jY���y)I6��Z�Q�I@/�����a�I��|w\Өf���DdtX�Ql�i���~�fd��5�,+=�}V~S�@P�G���#�#������2��ƪ���p�[��A3��]���s�i�S3�/�3g����6��W��={^7p+6�	*҅�<�2o������BE7�Ô�N(l﫭6�̋�������8�2/���Pƣ�M�j����i��$��,m*��Z@�P�4)Nz�
������I_q����9�Nʳл�~��~����k��t��.[c-KQ�h=K��ϟg�%y��_u�� ���S',�F6�y��2 ��U[U,x���/��`-�j���-]��_�k`Y3-���K<��'X$?�`��m�ubf̨e������[�����y��--�������TWW�,v�̙�aÆ�w��?|�pMSSǌ���K��;�t��^��뙛N�I���x_}o:�ľ����;7K��0G]�P�j�$�y�>���[�    IDAT���ysf�Y���O^�vՓ��|'��-����E/lٶ�������S��56�K��%˕�|�AXZ@��$|�R�`8�ǊI
�kIiY�z�����ω�E+�Y�,`@&�jt��J�w��9U��|>�U�1��Xl����$�~��T��磻���[���c�Jh�u �c���1/�"�Ţ���,���!L)g�1S��c5a��c�6ט^;�"�����Z��9�0D� �*�jMyy���#�����;����S�����q��[^���=�f�Y�\�|u���>W
��ݻ����%�;�A��u���(b���r>
�ٔ��:X��ϼf�PU��d����h�@�����|�ɺ�T{ �X�;`��>�گ���G�s^��~��=����}θX>��+��{������)��Ny�>�w����+�^�g���l�*ʫ��o�]M͍6^|��wK��>t��?,|��b��@�\���N]z�rϫ.-�������V�(�kX|����'M�9������\VZvd㦍['L��mJ픃�����GFF�?^�.Og�L]�>�w񧱱������t�ڶ��뺻�/O�����S1��f��<��uқ���>).ŗ�Py6����WQV�����ҋ������xi�٩�%�~���۷��4�S��Snn�M�ī,Uj:�F �2&-\	#�6F]`-����+_W��rY$FE��c<��Y،c#<Hޜ�������aluv��1'#��G�^�n	^��� �9F�#�����r�/�8���y/m~�+8��7�i�Le�D� 4,!���6��k��M�W��iӦ�󬨮2���?�B���/m����|kK-v�?sk:e�$C��R��  ܧ���x*@z�Ѧf@�í����_l�4�ק鈬V�w�nt��2w�ɓ�0��ݲU���>�E�Ǩhڮ�ZG��@j4-�g���ʚTic���īs>c�҇<�J�ٌ@�=ғL�1*y<F�3S"bid�y��@W9@��~���ǭh	���_�6��)�">|��y��V/�0f/xU��~�-u��e���~zoq��y�*�x���������_3��Al��/�}B�Z�^�t�)>�gβ�Q��f͞�4}������=��[����Gn�馆sV���m�u���mm�7tv����׷���uj&�9�V�)��)���e�
)rB�BP��(.��rv
�:��z���i��7u��w���~����-������={��lh���n�V�ާ!�CǇ��
��52��@� 9��B��P�X/�@^���>	7YȢ�u?�{@
�d�<��f(�D��1���RdA�r�{)��u�~v�ˣs�"HZ��^��]�/�VXc8�
Z���(���'-ZԬ)3%e�f"U�jl�v� �CyT)X�]�&�=�n8�TU�bӵx���x0�l��J��z���6�Cʻ�����~�U��W�CkKSlH�5��S�y��3/���	���/
��E�f�S���k��3f̲�Tr�����j�3s|�w����9)�����D`��y\�] ���վ��R�57�h�U�����H���`:`]�,� ��u�ڌ$v� d@��cm��_a��{(��c�:�(ݹ��#���r!��w�sڜHr�f�1f�<�?�g�eX�X�ths��<wSj���Ɔ8�s����YSb(����s��}W��Fl��62��'��]7aڄ�+���c����Aɮ]�j���omoo���em*�_d{7��%��:r���r���\wS ��:�bc�BE9BE�9}F�3{��׬��E�W���Q����GFF�^|e��#G����[Bssk���hNF#�UE(R�T�@%`�p2+�HL��F���6j���%��%���W�)eɯ~6�X�o��:�[a�3���`�$���j��De&-�����'�(���Ƒ�N*:|��o�S.��#(;ِ�Zaj���a+f�.�����j�N��j�>��揰�.\�<��(���(�"��kZ��\[VY�m큔 ~f�^��{�����z���sܽFwO��UUTZ-q�g��m�+t`s.�q-�~��Ϳ <g�oE�W�+t*)n|UQj������3��b`���l�Ȫ��b$�%��9j��v(�'B1Z҂��]���
s���
�����蓎e�sᔕA��T�?��ec�p�ͮ�o�D���G���kϿ�*̘5��ܳ��I��V�\�,�X�Uq+K�.S�L���#����}�]0.Cf��<�Z�|��'\(�o��ɹ-��w���*N���XE����R��w�=�~���/^v��,]�x�x��7-����;v,���������z{{���9��3D�mil^��]�]2�(rW}`v�P�Ve��[��nӽ�~�l��_k�Л���ܳ� �� z}c�}E� ���%����������Ӛ����MZ��!�|��%,��,l4��a�h)���_���V�-�	�m4�8�S�P]I��Oq�@*
���MYҮ��T��Q�广���^&�k�驪���������|�D�k] m�K�|p(�t/e��p+aZVf��A��W����Q�?�{�ЍeV)ɱ��Y_Q�`� 2���{Bii�%�
� L�#%2����-p�Z־y9V�<QNX#�A�We.��XwR����L!�
k�8���q<�r�Q���T�S�EE�����f����Y�BƏ5�8V^Sl��ܳ��w+��gMQ.��w���W�s׾ў���gR��G�]�����i{.�	�Coc��aH����ӿ��K�*s�uÆa�}�h0_ ���Q����v�	8r�˳�Cu9����$�{��+�X��.�0<��/�/��EX����K.�x�ĚI��R��.\�m������4?��W��^���������z{{.�D3)�m�������5V���}�fL #P�+G�wŧ��&O��㖛6��f8��_�W��Y��S��ݷ��X�t�V�X<m(<���ڡ�On~Ռ6I��E�"a�`.��A�J�VVzl�ܣ��l��Y�mI�ȩƆ\���&�eOo	DY� �L��_@��4A����z����\�ѿ'�5-JV���@,�@��BY �F,�z�k�l'�âf�}i���5_������:N�0�- d]YK �ݛ��&�W���4v�̽��53	��7�qP��wK�}��եK�V3֖�%�,W(@��3���\L ���A��Q�P�`ƜH��\��r�D�L�n_�銅P��6뱕����#�])p��`�C��h;每�k,�k?��y4<�Nu�ݕ���󒊀�+����2]��L)M�R
�����߇ys=h����.�,��?0j�9�����Ⴧ�ZD�s����1Cc %��J1�fLO=��)�'�æM���|������XD�<x�_������knO�2���:���*����݀:{15��?�~��))��e� Λ;g���ܹ|ɒ���ߝ�8k@�w���<x�Ϡ��_��פ� �p���c�����Ru!�@h�uߝ�_'�����.N
T�g�)�=ɱ��k&�%���dJ����G�!����2e������D�;��8҆ �sE�� {�Q��� 7�)�"0�I�
����PYU��&K���|�#nq6�ۛ�k�Fp���BY#/�o/t*�����^Ƴ�<��α��g����D����a]!���X��?�Os�6<�螑��˽���T�[����j�UW;v�̓��%@�1ѭK����?��=�Ϋ�=�Sq�T���b)`��'L�f"-ͭ�Y�Z ߔ�7�7���X�|__Š0V��/����������>��`��o�"ʹ�=��&���j�����r�������O�
D�F�A�8�o�����qCé��J�������7szm���v�m�iN�(�:thځ}��ώ�·x�:::M��~eCՄ�a0�O�.�ɪb����M�r�vڔp��%[/_��΅�窿M���}����<z����nhh�r�����|FKi�1�x��Kb�E�K��3 �q�p%kA��DBV��!	����>��7i�[�f1Š%,t�F��퍬�����s�{��E��H�.�N2�꘿aAk>J�bl��f����yX+���,S��.49�u1�~�Wز��X��c�?�
�����(eKt2/�]�������>V�w�r8���5�xD,��|����J�9�BeLCLwBI�y��%ʁ�~�)7�����U��{���+p��mĳ0��f-��%*�5��ÞDa�gF\�"��t3Sv�h���PQ?�5� Ld��D��$���(C����W�\i_�Rd4~�[ z�u�� (N����sX�g�}֞�)��z��}��~��Nցq-p�7����X��������X��"��˖.���7]�Go�l��[�O?��M�M����[�����l���u�3QV�m|�6>� ���iS��i�SHC|~���:w��wt��[��o��з�ص��������e=eZ���`R�V,[Q�x&~�,�&E^�����AO/ڱ�w���%:3߃��+��4�~�����.�\�P�	U���Y�\�KE�)_���{����/���yæ��3sT�悠�5i��6��|����ߌ�Nk�di����s)2]��t<�Vw������# W]x,fQ�^3=�m���"`��\�c��Z�X�r'n8潳�xFbN x(w�{(w��b���\�C���n����غ����@�y)3�&*���u�ĚJ!��8�۹�z��3G�Ce���X?>�B(p�{�(��Zk	�-�1�=��c��O�[��V.�c����ޙ�'%��[U��0K@�Z�-[r9�4_����`x�Gl/p�s�M7Y�j�>�n�cǎĠ��P���g���|%b�������5��J��m+�4���������u'�ٿ�����xuuw��������Z���0 �i���E�?�{�?//o�3��6��օ�
�GFF��l�y����"ܱ�)�*@w��8�C�!�hT�I�����(��Jz޺�왡A������!50h����	o�[/l�@����-p���M
ȱ�SVU��4��:`}��|��8 �}=p���N0���+bz�L��f�'M�`��0LL�R�:�Y
��lZ�56鷴7������sQ����<�N;���~#ˁ�Lt���v�ª��Q�b�n�2�9��ͫ˃��im�u��1� ���`�BƇ�|�;�rnE�']2�s���'+�q��Ϛi=XOco�l\�z�>���q_֚�WՋ�������\M�9s�0)�gi�&[���GD�9��^s�59�儂0\[JT�~ϜQ�`�����;�y>����ިNm9���f����������!�}���g
@{k[�Y�C�D7�Ͽ o4;�����Ym��}�ګ���{K��g��3������ߚ�Z�54��]�v{S��:����Z��0�xo�Z�2iAra횵��u�>��_�skg���#5��<���R%@�)�N�j0� !�Ρ�c>��
�=�\�+ #jY�q��P�T�V�]+N�Q��"�-�=��5�k�SA�,+O�F�F�3	�:�җ�H�0�l�&$���Y���s��̪��ļ�|[~�sm�r��h����N��d}�g|bC�a�+i���J��Pp״���>�Aj\K����ƜbWV�%W#_����cԻ���Q���gM�oN���u�ye����Uq��9{�,�B���0+|حU�K��yn�I5�9����7�A��$p���0��Gp�S�^� �zT��^�^�F h
O��GԳ�/�c���S��1"�>3�$�|8_s\�n��#��ܟ���������C��.a|3g�2
�{��^N�e��Uޖ����o��1�6����o7˾��[��ߙ��\���\\��	��߄	��a<.Z����t��-�8>�7������C��|�?=����Is�̜3�bwڬ�B�e��;�q&d4���M�6���k����K/�ٛ���1on�
�S�Ԝ�;v��:�~�|��������'��,9	W����u�!��|�Rzjwv�   ��,�Z@.?1 A�G>({�#���$�w,��"�z������ߐ�Y�1�O�?��{Y�� �&-D�:x{T���SsmOJ,n�ŅP�%���(0�rpY�y�|z����hk)%����r_9>mK��,��7�0߀��ȱ�v����ueSNρ� �[����Q`P?V�J��^t5+�r�xE�T��.��Z�,oc�yǲ��X
 ��`�27.��S���w����O�SVLQ��!6����b���Ѯ��76�A��3ȉ��	��Iv��$%����ܗ��*ך��{�׿�uc��T�k%n�}��w�o�۹9pܭ��jmHt>���ε`gl\�%F��������b�|��O\��q����s{�N޿��w::��Ø����R)���]!û�w�7Tܿ�4}���wm����;o<=�-z�g����:�tkK�	]��M-�
�VX�iR�R$�R6p���Vp:T�_�$�q]_���4z&����}���9�#��2?q�R�`I*�4x���Vʄ�퀖�S���Jϸ.����S6'�)(s�*06˻�̄���[�B�`���R��QY3���t4*ǻOשa��
b���t#�^W�Ĵcۘ+csK�A@K�݂%��|��ݭ��<ϵǥ����� ��q� �ro�z=�]k`�1Ls�	�=�H��'8�<?E��3�9�\����Y�q�eB�h	��k`L@��5n�js\oHAq����k��Y����X��Ζ�R����h_���z�0�?�-�) ��e��;�����6�~@ �L���Κ��:^;w���������hr����W^�� ���Ԉy�`�':���7J^�������/Bg{��Ńk�۷'��y ikr]y/�
cW��W]z��6���[$��/�X�����nCC�G���N�t��s��&鹦8�{<�Y�5�a�����}w��o~CW�� �Tc�mǎ�aK[�	@
@ǿ�כv*�ģ� ��*� E6{�� ^BO���uj4qO�xcS}x��Å-���~�T����U�R�8��g� K��u(%�����e�
��_��5&�A2�{�&�Zjnj	UՕVm�(P@��o���{i¯,�5v�P�o�;i�r�J�Y��<��3����*^2,n���*���g�eIٱ�r\	Y�ߦ�h�w+˸�қ6H�R�jlXc�y�U����OUX惕��F�T�c!|� �b+P|�^���ύ����D)��ȨCX��H �������pRy�G�r-�)��v��Wz!*AtkH�����n/���!U����Oֈ(s�Y�� ]��D�Y�C� �.6b����=�裹��:Ϝ1���u����g*$���O��O���a�Нms�� ���<1 }��K�ݰn��ޕ��=4���������:;�6��ʖ����e�&3F����y�����=od��k�ڴf�3�%{ۦzV�~��ɏ�8^�e �3t��v�I�ۓ�2���ˍB�Zp\q�`.��tY9��G��%pa(�◿�eXr�"�����B'��E�w��n��q)�GE�&A�c�As��|�N�ǚ�Yo�����#kE����9<���Y�l&�z�s�) ~*(
P)�*T�m��A,pf�.p�{0ݟZ�K�X*[o����sU�b��"ԡ��*0���t����trP����;�!��V�,QO[S�:>t��z��Ěc���sV�^m Q���=��@�@\��hn�@N�ɩ�ѱ3?,�y=@    IDATuO��)I��߸���ąfJK_�G�Ө`�U�h�%�b �Ɠu%�{b��꽎"C�r+�!7GAA�O?�C]��s��uQ����^`٣��_{����~�zGC}cرc�=1AI��[n����N�P4�,t:���-�"�������+��b��'�6�6~��ؽ����G��cCS�r�%y�QЛ�[m�d<�:������p����,\�����3^����G���'O5��8B��b,t��V�����1�΁�4�{Թ���O	b���ܰ|)E��Y�|����m������*��A�i�l��Țf��B��������1�5�)dRds���;�V��n�U�j��w�~��cO�+� 8Ƈ���>&�(T4�Q^QT�5X)���7�u�+uňl���|� 1u��ȯL� [�#�!��
um`�����"qT֮�O�8*V�d�nH��%��.�.kܓg�f%�' �b��}�=��]*\+	�b1�ֳ1k2ֽO�9��|�y���5&O��n�._w����{����������s/��|SHj�sL� =I�ˇNښ#挂��(1��y^��x� 4�X[�El�=�����R& Nk�J���>s@��4�@�3.�6m2�t��oX��a����F��x㍦P�Fh�X,�J�;֑mʺ �)�+@_�v��]���3�^�'�S+�w�ދ��?���u'�oݾ݌��i�j3��6�J{ii��5W_}�7mZ7�~9�'zV�����45�ܙtj�#8�RI��� ��������J��P4l���K-j(���u�YmX��P<���խ��n�`40�l��9�)�\2�ӗpT
�Y6�rH�������Z����VX����܋`+�'B��{��x���6�ph�@܊Ȍ���
�}P�Lk��!���xsEv[��o�i@���m�Qr6�XP��
(=;�l$�'D׳���ʥ�����
u��U�J�މmP��˱�9�G�,+���<d������,t��\(PN� ��^>t�ݻ���o�ŞE��+v�U����C�´�����s=�_K��?��}�
�_O�W�sD�a�+(����󈽸���<Ooy�bn����c\W�"���b�{�r�W��@: ]ŚHD�� ^�j�ב�(���]�m�E�ܥh1/ �� ��oظ��K���?�Z���ÍM������bq;eVͲ��׬t>�+�U-3�+���K��x��W]t���&.g�<�
���ٷ���}e[G�	lOO�	�t����a�w�P�5Z�t��E���-Z�z�
�����ᮻ�2��d8(_*��KJCk[s�f̲���v�52ZZ��[v��d�=s���,+Z.�Z-B��[]�R�^fVp��gFj�k�sM� s��j��f��J��1��|�Yd5p�M�1��K����α`�`5�cZ���M�W֣��5i��Fw��Q��?-�DEW�Lo @��>P���),�$�5ֱ"�Cձ�*k� D֜���eio.�^��k���Ɩ�]J�~�W��R��|��bb�_���|�W^��ސ�GSj�O�2)̝3=<�ԓV(�r�(�̥���:����r��C���y�BW�>����`�,��?���Ag]5_Y�t)��%�c�v�Y����Aɇ�\f:��\a�=���KM�Hu�%��`.�!:q����/��*R���p��MK�/_��,������
����������;B~��Jvvy\�- 5�YQ ��9�vZX��?��������;fHg诽�z][{�y]]ݡ��+��^@�,�XrT<�R�nn��%.��)�
�@�̊+��tk[G���:�:mS�6:?ňJ|��>򡳁�rŝ�<k��,�~���c��R�'(�bl��Y�4g��_��X�q�/p��&E%�|�1z���nd���\q������|�WQ��썶O���6���P��J�r������=
BA.�\�� �J��}����0�@�w�� ^�nƨ�U�����Xǟ=����f��B��-�m�n�3�3�)�=	��c^D�;��:�C��$��oa�֭�&M�2��{}Ѣ%F�S�����T�[�b�=ӽ���b\x�U����� �gM��E��W)�C[Rֆkci=z���=X>��)]�Q�̟����E�g�l��P@���O�8e�YP���Nk��9�)���ٳ-n��P��~�s������h�+����m�3g����kο�����1�r|�oj+�l�񋃇�=t�gФ�m�b�K��ZE�☈�ŋt\�ͫ�/�7���M���|�:U�v��u���sjg7��,t+�:8��b���7%7*O�L�,U]l�2���2� aE.���͛M� ��=���u:����P�.]З�54�}���Ƙ��{$�,����)�V@���j���{���_��.*,��C�n��7q�d�h��,z��c;�̼,�h8j*��xO�+�| �7��Ҫ1*�SҜ�66a�˷B�p]��R+(Y��������p8kݔ����(&|�.
Η�U�����H��])|r50��X�Dkz6
d�B{bϠ������H9P�t���:\וύˇY,tz��]{�eR�*��/+/]a1	}��y��ŋêU�c��m^5k�c���"���.�����P���ڜZ!��|{F�O���3~*�q��8�������\ce��Λ7/W�5�Ս���(
Ģ����"p_�������㫱L=�f�74��Xt՜��Z��F�b����>k֌�����ŋ�:C�5~�9������}�����K/b�S��ت(ce����*�:��Y3f�������n�q�J?�g{ƀ���Ru�������Y9߼�n�]��Y�~��(�a �Odp�ih��΋/��������+�[>0UT���� 8,G�f=�Ëңl����N'�Ȧle,�M���,�̂��h�H�.�[̃R�8��)o���PpfϚc������L��������W��EkҼ�c�� /��)(i������[2�̀5Z�
��`~V(�d1��o\~X�75��;)^��<������9+>��1ܟ����)����/�@0����A�>�Ϲ��yEgs>�Q��T���;�c6%.ߕM���9��НlӦ�Ͳ�'��NS�1����S�����V1�ʅ������+|�{��k�m�K�a�U`�\�2�.?���M�bn7�|����F�3�[,���{��Dse\���@�߱.�Gb-�&��|ۭaϾ�a���Ma���_���/qoшe�Ν��܃�e�&=���$4�49��΂S��w�L��e�%aB5n��0o����ٸp���g(��O;�W�ɧ���������l�f��'�O��>��F򶲼����TU�U+/m�f�u��+zg�p��{zz�<t���������v%_���Y�Y���ֱ���a2���｡��uA`V`����߰t����&t Pk�QQ�K�Uf�-R,G	j�z3C�hn��)���z%�������~�
(��P:��a�ZST�N���J�'cR��ÕYP)C��^��c���f��۸�;K��\q�������y��S^��=()+�ɺ0�$�U_�����0֮hb��
h��U8j'c�p�Ҍ�� _>w�]���z|�������c����d��I���o��jY/Q�:F���]ʆ�S��:�kб��_u�5�|f��?���l�E�ƛn_��_���~���{L���7�い�r��|��C��:�.@�>b�����h�BQ*��D��@8sm������;��nŞ����{�����/	?��aΜف@7��F��i��C]�0N����:ۺC]�Q��[ۚB���ƴ�Y���

�BueU�:m1-7\�i����;�Lt��u����=�flݳ��W�n� =�mC}����
�����RwM.���p��W��5��ҹ>�sq|g譭�Y���$ N���"U��=�@�T��<�A
��V~t	W�fY8�7�G\���5�l��taAk�M+4�,5h_��Q<���=D��[��W�l���UJS$6�r���a�1s�����u��0~��`�!���'{5��wCS�_��- Z�� yԺ��/��&Vט�&b� >�Z��ey�4�f��-���K��6r�E%���$��^�bG�MA�*�l�|ҹ���o/k�|�Ş�(����j�3Wh[�c�T��kM�4����6�B�;�3@(�Ir-9gt�sĊH1�j�� �B��I`ֺc=_�zy��g�51li�~�w� ��9��<�1k � ���'��&1V�wh}ѠǷm��x��v�$�?� �(����s}��~Eӯ�|mxꩧ>��@����X�ի��O?m@O��{\���0N����)����O�� ��<��`�wq�Yc�ӧ����ګ.�?�G��ޕ+���my��/�;pȺB;zܲz`(�Ms����c��L��^�����p�ڙ3g�ޕ��6N����c'�Q���}��"\G�
<�zȃu�9:U��"�y�y�`� �$������XN��fxl��Z��P���i��)����4�5����2P����B�˹"�<�%PUMS��0�v���&�sǂ��V����*�e=�k��Y#+
}� :��hb��d
��~�Uz��}�^��/:#z�k���n
��z�?�?>i�b�'��X貆��k,U:j�����
lK����v�P�,��?�v���E�vv���)�jJ�@/���u��.wEеrA��e��Lf1�qc�[�F�


)��a�&:�5���w6�7e����=���pϽ�e��=���X]i�#����XjO��G #�X`�я~�@��!
_U���ǘSr�
,������z���F�7ʻ�1�.+3���'�����n�cQA�h���P���uv�����Bi����U֙�b]*����)¬�3w=���}��(��/}�@}}}��/m����//a����R)�Oa-+!��$TU�[U����k�.]��90�w����ۗ�?����9����m`�e!@wk�_l�,ԬG⺵N�k%����Q�b���òe�BiE�������\�!����̄�ϥ-�t	(k��1Ϻ'��im]f��ə$�l�<�&|���L6�8Eq��f1'��bl -�����P>8�9�= .�����P�"��V�Ef��f՗[n=�
�˺���m��a�Ϲ2"�
d)�i�zcڠ(w���r��nY�O� ��Y��:2|�0P�x��|�ke5�]�cVq��I��`�q�Z�;�Ѹ���+�s-e/��E	�wY�&��tʘ&'��1�z��z�%����ؙ��H����0և� E�� ,ʟ��M�<y�Xʷ�]���&t8~}�=��H�P,X_|��t�Zg4�p��B>�uŪ�V!�H����6G�{���۷o��3䦫�籎(	'�N��d�u�t���n{z����L�2@�4��(��?�;^�����=�x�W?��/�w.KJ��RkG{�hq��H�,��8R[7�|��7o���3��{��3����뎟8������G1���U9�tYW�D���Ff�G�ˈJ �3Y�[�w�7�(�$���B6K4/�(Q�N @EZ@� �����V���� ��$��0~�~��-טv����҃��V��FAA�RA��rot���>��|��P� ��wZ�9ׂ�'�	k�v�N��r�l$�S�x�7@���3���5!�OMZ���D�<��	|� `�%��'>���Ql&�7�*�����-~�S��E���X<�ܹsl� q��ښ�j� �k����<���\�Z[��� P+>@��Al��{��������U@aC�_��{�����q���M.�ݝ����[�r!�8Zw�
�#|D
��� ڢ�y��*1m�X˪�Z`M+K��(����']��K�>y�2�4RAa`|(�կZ}�������;B�u����}��XTJ���N�j�:� ��cǳ�˕�o@�>c*
ʓ�ߵ�a����z]]��-��x�ɧ�YB!(�lcKsN�7�����*�WU����/k���;/���mz�,�[0�3�'�>|�ԉ��:�Е���*�̋m�:>�U���#1*��c�g�~|��ѽ����3#�6��@.K+�4����y�30��Tw�7� ��;onn�mN��xMv����P��ץ��v�Y>�U5���L�(���܏�"��N	�T�[1�,�ZLT:�x�2�������TU�� �����E�eG��?j�2�5��M��e��bG����X�貊E��25��<���^��hr�/ �?��c��������\�؋� �8��!��Y�X=�]�=��A�%�W���-e��Ӑ+�t1E :�"�@���9=�P(��������L4˔���?��4v�3�%*M6����i��\-x������Q��ϓ�wW{覛n�`6�n(�����~�#�տ�����	��_p����O��ɽ���s������\<ϓ F
����&�WWw{8~����Ԉ��,.5�X	�[�hѷ?t�]zd��%�+��s/��'����C�3{������!��)C��� L�XΟ?/�v���[�r���|�Џ9�'�O��ݽi�m݃��\D�X�N�䷆*��V���E�W�n�bt#��^9�� N�3;$/WJ0i�����?�<8��(�n)<��6�x^x���$X	!UY�,���B�0�-�"��'O�b�ˇn�6)�u��c���2�@�8��p6{9�yVR���*�W����VhA�3G���u��I+ZV)�u�a4�mԂ�ml#-�tΗū�
L��2П��v��;�(u��*�M����,�H()�3�^�e��-�� K�%�������Rlr�z�劖g��r�8Ȃ=�@OZ�j�BA  }ݺ����rמe��f����;���Fi�#G��5+$Z�D)��аu �Y����r����y��lr_*�}�s����W�cN�A���F�����Lx���w��]����9Jq�y��7�S��Tؿ���M�5y~q�������_<(w���{F>��u�-�B�b`_'A3�Ԫ��p�EK�����x�אUㇾ�W`��}3�m���^�3k[k��������c�f��ރ��'��o�n߼>//�s��?��8c@?u���'������+画wq��,P���C�C���xH�¥r�����/��*k������\����sY���\� ��:����BI�׊O��ϯ�3t���Ɔz:�ړJ����di#dɣD�U�L��% z�r�#��u-�Ht�ȇ��׈�T>b�UB�zA�"�9FAq抈�Rs�R�7>�nlG̳֚$-r����r�:%���oN��m����k�Ef��$��&+����_ey�h�w�r���������������)�Oy��y�e�'�{�eB�g�y��=*_���Ys�=��XkH�.*�7��Y��vY�9�A-\4=��eMi).#%�8�g���"[;Qٌ���js*p�:�=��s��/XC>�u�x&4V�KʞUv$�w�}�O>����%-(NM|���}C1�}�
�Y�zP� ���0J0-��(w���^�x����� ���Ua��K���o�����?�]��������!�=]�PV�x�A�������a���MW�Y�l�+�Ex�'rƀ^w��gO64�~[��E�' ]ֶ =Wtm�-:����
�/�?<bV���'M��N�c�����hf�]�OX�>�9)N�^�d�X;�ZBwgGhjn4��~�C��l-��������9@g��ُZ���䆏~p�-w(u��d ��&�~|�\��ѕ���    IDAT�7?dl�ɃJ��@� Zޜ���&(iY��؄%�G�u�)Rj1 MEH��\'�Q�^�<�,X`4-V��|a@DsDM���ٌ���4���IМ�ҙ~w+��Y�\����$��"�]>u��uP�:E\�}�����-�ªU�������J�D��j��+��"4�6��_~�
 ��(�`���gM;vl��]^|�e��T(p�R�>R��(���yuD
17���>�1��+��b��e\��k�ꫯ�.�����|�U�htGZ
*V:4<�O}ZZ�r�k��w� �4Lk����е�Ā�2SRhԜ�f��W�����ŷY��_�Z��_�~�O���6������zR�+LP3�ɓ'��ܸaß^���?:��qN���ẇ�>l���gA�V�W��xɓ�n/y��z�&����� ��KKsiFDgK���P� Y�@�K�<�V~գ��
���MMa �
Ǐ�.e<P �\X�n�O��UTs+�����`��G�;T$�o��iR�d�9�%q�T.E?bD�+
�~R.rty"�̢�Q�:ft]�ֺ�;>{��J/��J�A�R�r�[n��_iQ�='�����]{ I�[\CB���`?���������G,7������!E�kHP�)�9֢�]'��լvk+*&)ؼ t�5���c�������3̜9#d2Cĵ3f���w��{�@�w���W���ְs��ȑc���c��V����3��2.����%α�<�H���E�� 䀺�^ZR6n�h4:�p�]ik�����Yj!�ǜ{��q���>r�vEn�� :�e/%�1�w��֦f��%A�ca/Pⳬ�4̛?'�\��Ϋ7��/���
�8q��g?{v���_[�\�;�9�2n�Ms�M���;/��r����c�Ҽ����{b���$��<��-�mw��w���^�s+�b��nI@�s:T;TVO�r�#�����&@I��Un�Q�Rѷ,�]@gVJް�Ĺ6�ˎ������Z�,�_� �`�| �ʊ*K�Sq	�r���e3B'c��)
�Գ�`Av����U�ZR�����%��$(3�",�����f���9��Z;=0��o��������(5X� ���lh�U�c~�����\G���R1 ��iI!�I*'�}	��z��ڹON�������޲�Fxα��A��g�$�|�aI�6�r��1��,��yaɅ��=w�����	�6m�-'��:����S�M��OP����L�� H+������F3�u�3@����y������uޡ�9
˛9�� ϓ���3g��gZ�k���R�X'h�=�`��g>;�&��7��e���bORL9�Jq�-������9L�:�*ő�~�嫯ڸn��oZR���X��~�����_�S�a�<uʔO�'��@n����/}��K�o����﵇�?�r����9�|{g�:,t�XX�jY�Q� z��r�=��v�v)��ET4o���y�����o�1��=q���c}�Z@th�K������֖����Z�-�\�f���{�_Ueu���2p�q����*�q��w_���e͒�+b;�@�+�|�A>��m`EJ]�J�����ԙ�i�:Չ�r<��0YҜ� ?�#��X����2֣E������<r%X�i�k?8xty�
� S@��/�Y����P�'�A{E�b�>�â�X���I��ւp˨�"\�Js����r/���T�Ї?h ��o=lAd�^�)<�����c��n��Z4:�ӧO3����ͮ��0|/�c]����'>�\Fhw����T��)�Q|I��γ�e��,���Pz�~<�O���+_�Ks3P��ؑG}���+>tR�H{�|����:��s����2k��k�N�Ue��M�\�j��{���{k�lٱ�g?{���thlj2���-�������`���u�^���_����[+uf�=c@����w��,���3@W/ =i��g)@�Є��C���Z�m�q��,Yr�	c�[��� #�����
M���z�ޠ�-�<����f�twu���k����TXdDaV�{	ҡh�b�a��*ը�H}6)����i�>�)�S�Xb}�S��Dڕ`��fb�@��4s�����N��N�ӱ��B��%k@ *P3���I�Q�<G�7�fP�k&X�8 �.]���T'������ �F��,0I�3N�`��$�� ��s�k.��u�3&$+)�R�Z��Gګ�
��z�Z�G�pn��̐��&T��~����o��{����e��N|-^h��EE��5ݻ��)���
�hY]��`�w�6����"0P���^�D�[=��.�����,+��
�\CP�X����c{ |��aLc�����,�5z���#�<j�T}}�L�M�͐6'@oj�dcP�Y������)��a��Ya�ԉ��}��f�83�5~�;u�n)z���T�|�`Sss���ɹ��g����?wn����O���{�k���~ƀ�m뎃��􂎮���ny���p�r� �'}�Ў��OO�"���~&��� �%˖�ߙ����^a.g���yn�Ti�G����9y��}a���rg!�Z���u���o�0T������q���JP��"p��!��gbt7�9�y�L�����hb�rR�c#�{��h%8Y�z� ��gL���>W�_�S�����K�y��:y��Y��A�kN�(�X���K���wV=�4F��}*��W�m�>��q�\9�s��-w�@U�	bq�*!�˴��nŜ�3&�0?�g�w�jk���|�+f�ӭ���eghb�A���w�f�eKLy��w�����(˵PE��. (�+�d��+MQ �quPc��ȇ9b5c��T����܉?!
���43��,������mł� �����o}+l�|����'�,��YY|��\hl:z���������A����3��Y��o�k����moBF��.[�G}웯���C���;�a�`Vɳ���0��6\r��{���ΛZ�.[��|:g�۷�v��?=���#t�t[�`.:Y_c-t�,t���z���˖.h2:Z����
��"�r�-�;��P�z~�R���[Z����2Ou{��4V�Yt~�W�
t�B5Z{*͉��ռ�(�v�ЦF5&f�{�I���@N^�Ѿ41e�h��{��Y���I�ڑԃ���r�
�@�b�.Z��+ �Б�֨�uO�x�]`~���pKQ�%��G��q��J�Q���0Z	.��H��L��b���<G���(ڤ��q�3�
LAv�[�ODVa�@,t��Nc��.���{�o��׿�7VU��+_���X��,)��������o���5 E����3%���� ����V��o��K-��9Ůx֓�nK�,
�?n ������u���[{G��/Z���m�]r�{z�,���8+��X+�;�{ ��:��o8(��s?c��^������3j���}��M����K����+�˧���O��7��K���u����(�+��ZQ��箛W-_�����~�<#@)ܱs�ю����& x�~��ܪp�\D4WYPf]d,�ٻ�X���aꓧM0�L��_c��4УXlki�����^��T �PPk�\q"ҍ
��Bm4���b;�Ma�X���{@�><�������e�JI�B9YЋY�EX�.h9�w4�+k,��6a��b7�����+1ޜ՛�zG�0����8`�M�6Ũl�jP����Ӟ���=��+	¼thT���u�9���`�v�����K@
_}�Qܜ'&�^�W�D�+�<�~�_�Ѭ�X������]	�����՚slo��._��K�Z������p�-7�)S&�/����3���?y��)�?<t�Wo�R���z���:t���^!�.�k(TJ_�נ6;��yn��֬YcJ����P�'AhX�� >~K�,yw(������
qD�sΕ�_i�:V��T�����|u�K/�/{�������k107�Lh�K)�2g!fN��/����>pq^^�D�����ˮ��=�~����������-��uxk+�����**�bD���p��_�s��/;�w���Ћ���U���9�� @����%P�.V��@��Q��Y�~≆!�k�ʇ~7�F�?�\�`d-ϻ������;��5i劒�p�ҕ1����T9re!?x#�8c�O{0���%Y���5���E���ܱ�ՃO�Q.6@�ia�7�p��Кר1�R��b��	χ���@�\{wﲗI�qv�ֲ�ee����Z��F�W�-�C
�^XS�b����zK	`��#t3֥�4��-$���0w��>��GAa�+�B�=�K��t��=G�˥�.�؉�\�4���[l�ly)TUW�UWM��2 ��wvv��>u��PYYn����gϰF�:� k�wJ�`�G ��#��G	%����CԺJO�<��.��� ���،X���ͺ�{+�T����W7E��������Q��6�	��'BoO��V�7@�*�B�	�[��������z����+p�p{�?��{�N54Ωon�"3�Ǌ��>�7�@�2ڰa�·~�Kߊ����q��^�u��u�S�{z�Y@��`�Ղ�u��M�7�Q:����Dp\0�| P~&ȳnM�ﴢ�J4]���/CV�\R�HZ����MV��[��%MU	=�آ�-���|��q��\	p@��4V)	E��<�Pn���a�\+Ί��^�j�$n5Z0b����HP��8���~,;
���LV{	k_@��D�'AZi�c��@�c9Oύ�X�O�I�����NT��W[׬���{)v���8�{�zu�劲2��_��V��*�d�J/Ԣ��9�|�c|P�}��ߵ9�<� �����k�7F��۶�����n~�T ��ٌKY���w�ae[9�|r"��Ǹ�x�|��K�:�ϗ�L�25g�0w�io�=Oz���,�a<X��o_��� M��R��OKU2.��FBhl<:�A��|�}��=<�"L�8),Z����=x7������Ï>�}����L8q�ުv*�X�0���f����|��04��9s������+p��^�m��ǻ��&ttR��-�$�'A;�$�T�H�S�&���h)�M �W*�qm�G��pds(]�z螺QP���s���F�!ב*��Ï���B)�:n�f�v�EF�N�0�t6V�"	��@2��g�e%� ��T�H)6f����$���E�NT4� �
��/:ˀ��)l�\ ��J�Z�I�8��~��t�Z�c���b?d�s}��N�s�v&��q�!�^��� KR���k���y;[P�\lmrQ|�y����)�)�:��X���,��M��/�|.���6ۄ	��Y��4Y# ��6�x#-5��#ҭ�Ow�͗g��BU�5�/ؗěp���k.*��}��)��f(02�� @��ĸ.Zly�(���P_�͛7����X,�@�����µɯ�;q����Lhh8i�N0����8��?�dM,Yr���{��q���]���'_z����+
��N����\���7�i�1�y���ַ���777����K
��&TW��8iʑ��կ��T�VY��^]�3������u�����V��w�J@��-A=v�լE�X����U��Ty�S "ծ���i��F�`.kW�J@\( s���݁٭t�H��`@�O�0Ʉ���.� =�܂�R^&��I�2:�حl|��c��e|�Z���n�s-,+�Uc�\Ƅ���FKPp:�s�ŭh�쐟79V1����"�����4��I���8~i�Z�7y]�q�G�{i�
����I�/�&_����{��yV����^�{��fɒ,[�\�&7�{�!�$9��P���$�1B�i��ȸɲz/3����sgϫ�ز��5מ���e=k=��\r)��$axP���56���5b����@��ml��5�����/�_w}���~6oޚ0 ��u�ׇÇkB�;���;�g�s��+��{��;��j��
��l�ds6΁"�\��䉓�TzC!�ź��ɷ]����/�k�o/7�M�|�ki�u7y�����u���t����47����t9����&�5~��0�rX�;o�G�z˛��?T�{�Cx챧���#k>��ѕ zc��g�>�M��c�kP"o����@�Ť�ل�Ǖ5l؈�1��l�6y�W�M���ÇW�!��	zSSS�νU���J�[Z��3!��JӒ�p��6�>���o~gw��m�kE��h�X�󻄋Y������==^^ ����:eX�:��ط�{d�(�J~G(9��`�Ӈ�XJJ�,�wԨ1���������tYSn/��,�|O�*N���8e���tK^~Үn���\�Z��+�Kp���x�+;�.�IVjVR[]s$�������߽X���i����\boD��;��/��Sߟ14�����O|nb$�H���[.��i�������ڻ��ܱ��{e�����?���w����������c�=�����k�>g����ܹ;TU�c`�t��SP瞝���;��<b�����c>F �t2~�
�V�i�"7��D���޶������C��aMQF��sα�+U�<U����cF�M�߭\qNn8r�PhkjN�б�- �U��}
x>n�X�h��^x�����g=v֯�t�?����j��KTNR���H��"�n��&[��`�	UgF�xY��h`L��`F���l:e挧'����%�>��0'�X��m8���\�� �C�*�]�5��bUt�`]�2�[�o3�
QT����M��>׵�#0'�K����j���_ϭ^���L���{>����I:��F�a���qBYy�Y3�GD=�� 7?~����`8t~���PZ��;��z(�N� �c)�k��I����5-J��+n�J�@�HӒ�hv���Y͙,\�������"����$^ _Y�R�2��q���(w��c2TZ4fbeC�Ak#S)$(��3qo�z����i��M{��-�0���z����p�[�lV�Ï<h�;����~C��׿�Щ���� ����0q�)^((�v�
���i@W?xy�r Ԁ,%]�'�w�}��z����+ ����7��@��e�p����< ��3���/_n�;׃9�Z��q-J����z���t0JJk#q5��5\���<�Ѓ7�pN��Y�|��+�\r���¼�3�]��%?���G�j-^։�er}ЙH `A���O}�S�d�#
f�Ә?�O<cEA�0��Ə	sO����y�>r����>�	z*�*~�ƪ�������f"���z�C�-6�� YS�7n0
�D��z�OHu��*�u�ۂ���b����_��ߑ`�nJH���3}��aĨ�a��)v�P�Ny��E��/�k߷{��ny �����T4���nO�8y�W����;��-�ʟ@�:@���i��q	Z?�c�8���IA�Z��[�����b��:�#��m
�c���e�����;cJ��q
*G^�X��,tW ܵ�.Œ��C�r��9z��`X��E
���
4:T���������6�/ist��ZX�ܫ��x��n0*��b��p%�;ߧ�9焝�"/�kֳh�������x�3��mc�t�R�gP�����أ����XId�h=X�|/��M���� �7P�����oʅ����)�&���7w�������ó�R��Ç����\�?п``p`lj0�$;+�������y�� }YQ����Һ,��W�ھ}��Çl��}�mܼ��2O���R�WW^yux�{�kk�������XՄ�u(]4a��M�^|����<}�_�vڜ��V�9�f�    IDAT!@oH�ʫ6m������ohL7e������B�C���)��&��w�O?ee2ye��c�E� $KI��9����U�a`���H�p�P�6)�E]'f�}Q�����PVV��F�F�J+*-�IV� ����ۀ��ã�)�ɫ������E��*n0 X�D|=�O�[�� ��%*0��t��b*>s�2�zY�r	�V������5��pc ���}�<~��H��5�Fk��S��[w��?�rEK�~�C�}���a=H[�Jiپ^t�^����nE���(/9R����H�	+��r�f.^r�)e�
����\s(s��9�Z�]9�3e �FL����	�#�H����	�}*8�rX���������mϯ�U��m�tp<��3�&@�"N�8���>7���.���&<���IZ%ύ�b�>qr參VN�={��ON��p#�А*ol��@ck�;��򦨥4�7��2�0W%E%8M�����=0a��{*+����C=�̋�������,AA~��_�^EIE�D��!Bű����b���T2�*��Z`(�nĹ�4��e�ʌ�KQC�=�fg�v�x���Y�|�?M�4��*b�� ����bOÚ���2|袐c@��0 ē,@�ӥ���ItQފp�1m*��.a>�N��B��K]V���A��!C�E!kM�'�]�h~ai(��#G�	�ǎ	#G�70W3�5��˫�utwX����6/�����Ciq��u��� C��6���$���~�����<b=S����w��e)�/׹Ee��/ ֜�"�t�dν�wl��������L��������=�,s�ڴ�����|��cE�
� ��I?������ �tR� ��s�z��-�B�g~�k���:"izBPQ�*ւۆuA ?�8pX� A���{o����c��]�:��4:J���ߟs���~�!7ˣ��*�;g._�����}̝;�*ϩ��NS.�a��/��T���ٟt���ea��I�W\z��)S�4�����={^|�衏��u,�)�9v�'�g�R�, ����>bİ�M�����a���֬�����T�C��_ܸ�Ά��Q�|�V�
?�ُ�<(�*�d� �4��!\�(�ơ`�L�o{�Бǔ�����^��̍</|El���w+�u��)�^pފ�Zu��B�NP�����Օ����S�S�}�.�E��ꉭG�d��ߖ��},t&�I��_��%�%��� ��<��Y�i�"��(�[�e���b�3���"T�4@5ft>r��xx}ɡ�VW7�yݡ�~W�﷔&|�t�:PUm)v�gϲ�������h�mZ;CEq�1������:��>S�-������`���+�Lk]��)����
���ֱ����*�#��%����T{Q/�F���8M�'Q�V��|��Z��jXr��r'1R�{7�t�Y�{���]v��]�����O��6��>|4�}��f͢d ���k0@'���45�)�eP�&�����'xPŷ�� Hz��PH��m�&���X8jyjt{VVVQ�͛~x�1��DMz���o
_��W���G�e��ɞǕ ��50����~��`���F9���y��L�4y���o�����E�O��0#�i��?�>p�c�-� +,"���Z���yW���j`�C��(wq<v�ضSf�����h�O<u���??��]�12V���m�ֱЩ�h�'���=���w�ò?8�����N��e�{0i�5�����1�Y�T9�=����s?6k֬c��o��y�7r����:���
Bs��-tE�g��V]o�p��'�y��,`Y������s�>t�'��$N�Y��R֩(k�K!���;[q�G���r�m��t�����8%n��ߟ��%ehi�J;��}�,$����� pbճ��a(���!ˋ�� ������&�OZߍA[n�L��x�.�8=?=S�Z�R�b����
	�#�K�IZ�HB=[�Xp�s.�!��M�J��c=V��<���3�y�zR�^���mo{��WsKc8��e�{��cux��5�g�z���\+s�@UX�x�	% ���|�<�� f�h�4�#��I!Ch���]���_�g�3VzP�茆BD�:��X����o{gؾ}�1U(�@�Ϟh�K.��b�-���r��Q�fĚe�e����z�ڱ��Iˉʾ��M�����޾앋��G�&F`��=�l޺�C5��ɚE���xa+��`nm_%Əf���a?�$0B�\rYx����֭[-����w�?&�}��ӰmۖPW� �WG���rͳ�P�(�T)d�[�nqA��a>=X��Ǝ�?�i2!���^#D���@��ٳg������<㌅{����kt|�e�Q��j�3��u&������xP���=k�.n��� ��`�����&<�7�lg���ȓR��ѐ�(k1Y�,&=���3��&���|��P9lx�6<��7 (.�͠jY�9ٳ��ܟB��2�:�Vm-��k1:)GXs�͗����˶`+S@�"8����>���9�,t�o��Ȥ�c���t�˽�3�x��sI	������t"y�sF+3�� �]�bM���K���@o&��=��`��*@��`���?�^}�	��{v��+ϵ����?���D�k_O_X�p������閨������b�B���}}�?G���%k�R^n{��n1�B&�g���΋��� ])?�����]o%k�?�;��~A��8���e{>S������ :�_���m�;Q�P�6�y�W�G����3�������%�N��Տ����E/�{��[�o]{�m3'(e�uǏ+���іr��¨�mpb�-�����wZ�l���.��8pf��d�^���U��$b�Թ��|�_�B���CqIa�O����<�W��N�K��c��h�3F��}����ҭ�]�������'^�(�1�qB����<l׾j,��ְЭ�w�
��(_���<N��g���g�q�M~�.@O[�	�+(.;��b�,s������� �)jY������JȤ�t��?��������PZRr�]`��P3PO �J� �y�6~y�9���1�[�\طg�U�**vE�+oyw���<�g���P�_�X���+�և)(�S�$a��q�OV_�1Hj��yt��܏����Z�?�| R�b���;�%�d�J
��
�k�D���it)H��9oQ^^�ꪷ���/����o�������c���Ͽ�VDA��i�-����+��[�:,%����#���_r�%v��:��qRB4���.k�B���c-1�s��,Z���vb h�E�VSy�0�ba�*�ku�ָtr�cAq��Q�ϓ�ϙ����|Ӈ����]�ե��nz�[�l^���m��#X�qU��eo��y� :�����1̈́�.����a-������:=��M����g��h�zX�(�|�A	�=��ؔ�����yɊ�bwK�&m�����N)���VTPl{�s�7��D�^p�ʏ��o�����8!@oii�c�~,��؇S��g��K�eD�kr t�HIS;��n�9�;�Q��,�ď���b�R�w�\�>�Z՛�Z5X���F,�$$�hd��4�(*.%����<�������\`~D���XX<SAQq���	�Y�a����O=ƌa����X��yٮ�j����J�`�hk�
t�%��2����	h�4-��nu����@) �gF�� ��؂�7�>�2�ү�_V��W�k�z>݇�*�	��ƌ� Ae�)*��=P)���,���,����+��=�6�kim
��fT��%K-��Ӄ��-;� ���8<��S�HP\cs��O���Q;Y���3zIV\B����)�$�=�ƒ�}n·�ϨO��<��/�42���J�kQ_[[/^~�ӟ��2�c�Y"ŠxP����j�b�*+;�.�3~т����/�?�������o��g�<��TK�li7k��a�&�o�WTT�ȱ[G�	���Yw�E��n��"hR}#Ȳ ��=�z$���]֯�`�9�qnhj�\K�����������5���g���̥��(�޾����r�oֽuϬ�0'�9J���n�����ީ�&��G?���]���={����š��rw�܇B_�z,L(�l�+�w(�;�.zS���Mi�JZY�~�������6%b\]|< �� ]�&��V���S�ܿ���e4��ι�¢�WTZ�X �%V�PO/���hQ>�M�CӔ���g���9�9ܚ�����#���l��qM{��P�hP�S��O�q=�NM��AbEE`��(��� =��9Nq��̿�z��8���6������JyZ�֗����c
�|P�t����!ⴵ4X����]}M�1crhim���]���\c�����+�t��5����c`rt]�����O����Q<�y�~���c��`��%��(�c�쩧�K�f�餶����9r�]��5��~rs��{�uk�kp �߿ׄ,kV�����Ū3jdX�d�;V]���5A��x��y���v��3����<t�)w�?b/�M��F���B޷m�l}���Ya��~���i����<s��F��|��ww:�r�?{�ºu��9�u��ͺ��A6S9��
[�я~4����v�`O{g��U/�u��Q�'������w��+ʅi7��)��V���k)--�}Յ+��]����{�W746��76h��r�$y(a������L躵덎!�Q@%+��'��3�fu>Y�D��w��-t��Ꙍ�����M��z	R���,t4?��B��]M-��r�����d�M�}��a��a�3/.(4@��~<�Ia�5�&@O�+e �E�K9�bS���ӊN���߉�<�����XI�5����6m�
L��xb��X!��o�5�r� b�7�wG��H�F���'y�P��7�)�Y�_/��w���oyyY����J�B-��C�v���z[/�A=�'�V~puZ�ٕ
��(-�1�O9�	@��Z��+m�L(%��5�O�=�\۟��&��Y3��m��l�n��La$P�X�twC shΜ�U�-�tO 0�*p��c�� ������0n��pɪUg/^���%!��z������g�y�3��,T��02�?b>`� �#�Y�;����Ÿ���b��?Pz{�BIYy���~>lܲ��IcC�Y��m��_��&ﺺ;���;�j�(�P�RbY���ZU�������owo_��S�����-oyKXt�;�t_V�a��v��(#�����	&C�E�&LߔI��3s��痟vZ�}-�0��޽���������@g@�'�Q'9��<�KFF�/��8��-�]p�+�t ����	DL�4=�c�4NY���L�J+#�n�b&��%���[�u��J�U�]`n�N)6J�;F��,d[�_*µ�6��gB0Z���,;����xF܇�m������.�=VL��C���-��]J���,�������x4���=�JC|>���b��+�M�w�an*�����Xy݂�t���y�B o���bcc��� ��^O���$�s��̀���?
�������ޖ��� s��a�ڵfm������5�s��O.Pg=�P�X_z�ke5�=�<V���̳��\�2�������,�o�b�|��1�h�����K����>(���!{e%�q��YY��&E��0���F^���S,���.��M[�Y�}��̕W��M��ܱ�-Zh��#����K����ϟƍ%-���BXִ@�9t4L�4%\���P]�>@���`��n�:Z�C��}�!�d�7]��0���(0�r����ܗ�+VXL����~S(�%���%~�5�X<
��]{�$����-�%��WF���&�17���q����N����9�����.��F\#'��c��74�5�v������L@�V !jT[�W����EUWՄy��Y�^�hw��*����D0�h��Ā[�bb� "��=�I��CtPv���鴩SCy����W^��JP�����Tسwwع}��� (,'\�OlA^n�;�[B��߮�	��[h��5O|.�Gsû,w�b����z��^2���F�0+R�{�)k@��_��n���w7Cp�P�
�4- 1��/4�T�RN�)����Qg���O?#���Da(e^|�����uW�Ń����@R���P�?��C��y�;�I�E��G��o���0P�x�����<t�S����5"ֱNH�!����4	��β4:*�d�l����̷�X��@U/'�:Z[ByE����T3��X��SRG�	�7_{��N7n\�Q�!�S���K�y���ջª�S����6����`�
�m�ƍ�9w��E���e�����UՄSO]�{���~������v��ڛ���`o �i����ea�����*#.�/f��'(����7���FY�իW���K��%N�=�W��A���Js���t���fp%��L��0�:u�sӦM�g���}g����o��sB�Nd��������+�����B��'kO�[�
�M������� =���Bs�5�[N"�P,PH]�I���t��(�p���޻:\;���йk�Z�A#D3[4{�7S��U��,I��(���b��5 G�Z�դ;����|o%�� (77t���Ҳ4��琖ylTr�<��5e(��1�!%&f1���3��c2A�x�� ]`��P�AqX��4�,/:$K\�6�(`����x�,��ڴ&m\�R��q/ �	��Q���\=�W�%i�6#*���_zh�Y��^�YV�8�ғ�����K��ypY�	� ɵH�%�F�H2�P�������r� :�{Q�:�,c�~��5����_~���[���]�뮳�G�N�1_f�<���-mi��؝���G��0v�r&da�ŰX���T =��رc�.Y�zδiY^����6�v����O?�z0�c날4��;��0��N�a
و�
+|��M��,pE���u��Es � �YB�Kj0�45XJ.�{O_�2uF8���v>�L@�+����.V ��;���ۊ5���op[8t�΁�G9P�,���&ss��j���z�s�h����I3)�3آ�65{�SQQ��ӿu��|i�g��Mhr�t��oܸ����nD&�.���+��$0cJW��L��\0_]�|�Х����B�%�&@@��liet~���wd����w��>���c@W V�iIt%B9?/i�Z��;�`'�r���9�vg�SQ� 󽓷��Z�8�&�����N��庆�RH4n�{6i�<�b�|q^���:�R���Lk[׋=헲�cD����s�F�S�ul���/��|�x}��K1B<����<=R� ����{i@O�͜1-,Z|��P��]�d�o�[a��j���	�-���A_�җ�TW�S>'��0����<kB�	n��d��c�$V��z�-Z���+�ph>W�^8s��v/|� T�t��������m㠦<<��
�dg�#G��$���O_�����#��)S���֛N��-K}��}՛7�[�nZ^~q�m�O)� ����Y3�~@OG��c�:�Ho�\}�#?r�!lڲ5̛wj8x�H��o�̏��S�-t<�h��RHM����p�E������4�NK䚘!�J/Y?�яL	���[Ö-[,������y�=�\�q+���m})�%�\�O@>�(c��*�m�N��q�c����^�쌯\w�[��ܹs~[S|��^�����֎j�yED�0��[�:�g�u!kaF6�
�L�#������?�}�,4;����؃��s�V�( �?�ǀ.��(ߨ�k�P<]���^�׭=��Z�    IDATr�#T;��}6��܋�j�*�Y�7�0�O���Kܑ4�.*6~N~�)x�+D�kl�g.TSR�ң��X�8�w��1�Ǿ`����+��n��@�����u�Rb л{:m|��	�_�r��(/7�r�;,U�5��!�htR���y���߷��,�g�}6<���T���X�Rg=`���� ����s^RZ�1�ǻr�0�_W[o`-k���G��|Y�җ���G�l먖���X�T ֪(��p/��G��w��t: ����Q����G��s��{�Uo^��v'��#���xꦭ{6l޺%{0�Z�����묿��F�"8{֬0v��Pw�p�暷%I��n�(4���P����1kE�����VH����#���!���PTXl�s��������+�]�뉽�z;v��t��m�[�z�(H��D�������C��5u!.
_~����"�=&�Y++��Gw�ζ�p�pM(.(�q�e���w߽����q����aæ}G���V�]@ӽ��:���2���N�D�C,t��Z��
��~@�3Q��]��I��)"6,�-tYpr@��e�Rw��=d{-k���P
T�fB��\O�n�\�Ԑ���ʢ��H�7��K�W)�
ѳ1n1g.h)DlD�p�~<]�2�se�?����c@ϴ8E�q<T���k�C��[�[1����u����n�p:�;�inn}頸����5hY	,Q��ֱ~���#�8?�����JGa�|�Tm����9���|+�]T���Q;ڳ=4v�]~Ex��Gm/�KW��_|a8mႰa�z�W6�<8pȔ	� �1�����2s�X���aP/�q�;��Iw:%��,+)��?vL8m��?��╟=	���8t�����ޮ=��@*'�5ԛ�s�B�X_�:k��ȑ�Cw{{8���BQa����/ S-X�S���	�>�6�wv�#�kC]Cs��������J|ѽa̘�d9s�)�����aĚ��f��4^{�P��At}{g��q'׏"�e)�N� ��Y,��r���a��f�Z��bx�T(�ɱ�Jd|�X͞=���_u���=���h)���M�� ���c+XSڲ���-����P<���(iGN�;�C���DAq���9�Ԣ�E�Ě���J'�G�.0�i?l�w!�_\�� ��B��9'��8��s#�Y��m5�s�����,|��[bx�D	���p����Lׂ�^�\��k�X_̋|��[�1Ӣs�c��L:^�R�Ws����33\X��zH��[�k}��#�C��Ջ�]�ٴ������7J빸8/����be��njm��qŘ��
XP�����A��b���5����P���)�[�_����F;���Ʋa�,_~f8��塿�A�SkF�c��EI�:�7� -+)J+�h�Z�\V���	�Ɔ�˖�:�3����ɫ��w��qӇ���
��¡#���,�ت���A������.��<���B�)�2�H{{��Á��Z���C�`�#N�-ͧT�K22���3�iј��,^
����^��:���0���<�l�::�n%��ʽ�w�k`��c����ZD�{�*�(�xH���&�C�Y���&���xp��0�{��&7��/�������q�oj՝�ss/��~w}C㌶�n���nk>Cik�Lz����Lz~3�h?O=�T��n����Н���c@�F�'���=J�R��#��@�V#������:� f@��Hq@��'�H���%�wq���]��R��k<�-�f�n�s��@+�p���u����4& v����$�y&�-�H`��rK(�A�\Jk�j�A����Rv�䩳���<�:?�r�y�|  &��+��2��H֑,~����5��@W�`D�Y����6�P��{���,I!�kJ�o-Q�*���P<��~�-7����wB����nW̠���k_�H���4��ʟx�]w��C���s\��k��x�b[�P���s:`�j~A��CYJp�1�((R�a�<��v�<XF�nI�$p�{���ܱ�gN��[u�������X~S��w�:7n���/l� �������~���
�o�i�:q�ذl�顫���ҭ�^�iv��+_��16���3��-��k ��<��c"V�`�8q�[VZ�/_nk�=$%@rIl�5w�7��N�m ��ެ}�my��瑲"�Ts�sY�����;`q4�k!�ģ�� t���C����b����%H�=c���9��knlӧO��g��'Wg���k~�0������u���[�:Ӏ.+.�%���L�� Pap�/6Ҩ�LzL���k�ЙD�`�:����t_�c|��NzEҝLT���@)������)*����3�9ϡC�}�΢�s�����|b@��L��B!SL�%�Dkǀn�a$�EKkd���)u#����JA���<�LE*>N��5`k��Qq����FvK=�ce!��,tcPXiɸ�3'���1$��2���_�ν١?����BSK�	#�ɿ��o�>|��U5<�"��.��, Y�`�Cq�am$dEbq�V>�8��$���+n�쨽��6 ����u�}p}�(��ij��&����k̵>�?8�� ��ԙ3�5\r�3�M���I��5��7��ׯ߼�ٵ/,���	ݽ�����d�G�Kp��hΛs��'*
�;�/,/<dYS*6�sk_�jo�:VU{�z]Cc:U���������Ҕ�8y�(;� ��� ֛�ܥ4*0��1���I�Ē�;`�`*���`�L��}�y [>�a?�K��R7ȭ巳f�?��L��A���5���QV��=@�\�Y�ƚpt��¢�����ߴdɬ_k��	�ƍ�7���/���2�-�U[k�oe�j��(pU�	���А|����HW�K�3�/ʝkK�g�J�M���.�>�[�ݷ�.(�����5�ޓ��h�$�BV�(wiyq-��
�3��%�5>Z�'�q�6���K�� 8��u�3?ֳ��s;��e���C���֘i�ĊE샏�CV3����q̥@L]���������-�+��IjD'�dtkz9���0�z����9������p�-7��~��F�fƌg
O�������_��_L i���V�㌟\��:��<[�r�{`�zhOiΉA(�'=�e�ˍC�Vkr��k
��hs�}�rFAc�y�<ž���ﴧ�/����S@�M����޹��r@7�n��=O<��t��~���@�s��G	���	sN�i��g���n�Cv���
�=�xX�����Bg��9��A`[ss������PP��ee�X�k>��Z�Z�X�Y�úVN|&�&����#�=��Kh�� nsCZ�n����X��tP���4�v%�E���+��V�����E	�ʜT*�[�`�z(ޒ����`���J�J7����oZ�j�_�r;a@߼y�c�uu�64��l��|�/��i�L�g�	��M4�(a��������U����^/��I�ںf&�H��E��4!4�ApM��xzB�S���{�r"4E�Z�[�10�B[���G�$�� r��w-^�p�sQ��xVY����ФQD  6P��Pp�b#��+0�wb��>�X�o���/�t}��fLĒ֢���J�b�W��.@L%�A�+�#ʝ�R���?��.+�D�5����������=�����l>�͛�����nkI�W��8eE#pT>�{����N�u�+
Ę"��.͏�(�g���W�4�J�T��A��:b%�&��V�P�[�;�Ts_���
z�wܥPY^&M��O����n���_� ;y�W6�T*gݺUk{rk���� �`����ƌa��g�c���y&���?	����u7\z���+�,k�B.�'��[L��G�ڛ��I�3v�׃������+W�:V�,s�J̛����>��A��%�rTG?�E�~W\�E��֥�xV�U��{]�s�|r#c�%4�\L���F�����w��.�A=r�0�C�s��7�|���ye3��:a@߲eۃGkk/�U�.�L�D��i�2�v��R0`��)������&��[�ݝ	�ǣ��L���Z��,�t&�(w�l���=�@�Hw-�����3�]����L��-w��������������(_��e�10�"��=;ۀ@T]�;�;
��d@b�Dϙ9z	2�����$1��o�`B��N�|Ċ��K̍��!Y���4���;�Xm�h�P�����r���~���c>dVa>�7h@������3���[,�+���ZCy.�cL:�&0MV�l��95fv㉻]���8,���ѝPeor�LT:L
��墵k��dM���1Ķ������UV��>w֬�]y�[��Չ��G��#�J��֮۰���[PTZۻm})�\�l�r� Q��Z�ޮ;z���'�}�C���������J[[�dZO�ױH�="����m��}ݖ���w:k�W�b۴ސ/�\Vܛ�H�y������������l�����s�{ᮍ\c�ɋ�rO�D�&�?���:^�p5�|>��ҞE���a�]�z��W�Z������m۶��׽�� 0)��1�! -/@x����)�-]�Jq���V��BM����_"Խle�u�q
�S�$����8"��'/���+��KODB��V�|=
L�V��1�� ��ES�i0���-���g���D��~b�<�x�j�u,��̻��s����u?h��(B����X��d�>���6��qS�4��5j�k�i�xLe�j��z��|1��}j�s
U�r�}��h��bK���D�G��?4����φ��Z���Y�&̟{�m�{������a��*�s�X�X�1#D:��v���J딥o�g�`���*��k0O�'sSVVb�Cm&��l�f1�K.���8A���� Sg�#0��0�
-b��s�ZvފϽ����^�P�s�������Ċ�21��ٓ(|(��!?��c��Əc��o�����d��C�kj��I�mo�ҟ�D������y��������j+PĈ5�<�7ٝT�cmI���!`����~��w�k!o'��#�(�\���cE<`�Ӑ%�c"��������> �]��@�Ĉ}�b������������Լ�֝���\q��g��}Nзl����G��SAq�L��Jq�����'��oD�O�6ӛ�$�G$P��T��#��e��R��(�N@��Ԅ�`.E��#}(�q(��=7�)v�rϣ�ڱ�0Y`��	f���}a���wD�s?��i�:N����w6ԏ
Y��X�	��ʊW>��R����=��W����SMg��(����K���->&V�,P�Pv|�{��TT*�HA���=�o�/������3&
�;n�;�OZ�I��m��1ll�]p��oc}�	��/��$Q�0PS'M��my������|ꀵӖ��Θr(�ЌX�����,���-g����b/N#ˇ:��+�E� H��� ��jĈQ�?�85���/i����L�c;ԢW���l=�
���S��~��̞=�����ɣ_����]�����?�����{^�����{�����YY��	n�o00��˳@��}�k�o��o��%K�bG	e��ܹ�}�	�[k������o��`o�:yJ()(�ʠ��Yo�����?-��?��O�ŶXo(��e�G��ڝ^�^���mYR�˞���
�I>��B�H�e,�Ҹ��
�E��)˔����O6��܈��m6�x�X��������⟾��K�>����k�_����#G>���::�
�(p� =�b�Ad�;���鳜"�K���1���\@�@"�*��7��2�R�>v �i&Aq�ńRA�$����lBi�ɥ2����,@|��A�t��AW���lȇ)z�1�˱����J�
�/�R#� ��"�/5��\l��/`Zk�z"�+���~lYǛ*��z�F��xt;ǨN��+��� ]��f\KT=Y	�� �/�rŌ���_�o�0EeP��[�����o|7�T�O��q(w�z S(w�����Ξ�:��U�x���[ƚ�C�G�O��HY)N��
��C�`ۻ��&n
֬�{�ωB�?����D)vewH���P}[�F���}���<�x��J��aҤ����{�}��%�N���G���e���{w�6l�5U���	�K@S3��@����Q�=~v����������y����r��I�d@w��\����֎�4�s���"S�;�:þ�UF�� bQ�Xrm�_l���X�X�&x�b�S��'L���TY jwg����su#4�Z.�~���C4�؀J�Q��o�bqQV�9�܂�P�[`��~by
��u��_ZTlr���Ԛ���5��u��Y�<g�5�N�w����C��~��o�bt]�*W�������4��P�8�:B͋�G������~�L�L@�B@�r���!e�'7�S4���b�[���e}�� )(���V����q#���b�pB��@] ��J	S�a)2J�҂���9gE���+m��|ݞ�ݡT��8N� ��g�1ϴ��ٴC�S˸������AV�'vhܥ�����)�ж*�S�/�lH�`δae=��q����),���DY�;�Tg/���ֶ7���y���;�t�a򔉡�0;|�?��kj�{���W_m)�4���@#A�YYa�%a�̙���/<���֬B��Y�N�t:%,���pwGg8p�@hn�W��r{�֑���~b��y�O�����ʵ@9\�P%B�K���9��q�Ǆ%����������x�2���뭭�#�lٳ���EEqYyhk��3�P¼1 �a,r�!������/���_�z���73�n�ᦰm�.�׬O��XvD���T(n�	͍�������p�����^�:��u?X�C�@��.
S�L�FC�=z�:�=
�!�e���!y��*'��a�j�K������ㅙR�\������Šw��g���)?/���Z5O^z�f5jL�%|��A(�{?���}]J"�0��ݻ�֚C�JW4�;���N ]5��B����E��z�@�� �A4� ]BY�v_|Χү*G+`�A9�̤	fjj|?��% ��@p
�:�����p�ۚߩfϐT�3Z7'�
-��3=SC�+�N�6^t�]�i��d�8R�D��;��X�Ѩվ����v-�<�&8CQ̱��oK��73>[Qg|++z��Y��xq^ kS4y�^����smT�����t*Y��_��ƌЦX�x*䆎����.�,�52�]�.,]zz������a�O�0�Y:���g�>���Y�-�O�:T"�^�����K,~�^Ul���'k`��k��;�y��@��+Hk��d��'�ϫ�*;ϣ������,�T�)v(6�/ED��u�N�X�K�-Y��ך�{�¯��9�6zϞ��z��������Bw��j���]|�X�a@?Əg�K��������z�� � �R�X�)g`�������FIQ�lݽ^;��Ys�F��k���]� 2����d�g��~���~�;���^E���`c��|���u���p�I��X�[�X��l���\homMr�=8WYY����W�`L��a���a��Q�<MM���zXy��7�����k��������y���� �B��q@7+�jc�!�8���z��� �����q���܋R��=Y.�W�$k�{�w������C�
�y'4~��AJu8�[�ƑCi��M&z<�/i�z7 ��>�zR1�I�^QVn��(�k�4���	i��gSu;Ω�Sr"j<��=gni�F�E#$0b�)�?}O�#�'�D��|�n�آ��bm[s+��ub@SCP�8���4O?I
��L@���3�M50���yĀ�R�D�"9�m��i�
@���K��[yyE�+��z��AʗRθ���h�	w    IDAT���j�휤�0&�=�3����G�򴦵>l�^ڧi:1)<������1��ɱ��{0V��LEI�>e�����[^��:���gjk���رm�#�|��u������u%�� tw��y���[O���m^?����iӦ��3	��8W*�{߀���9k煾h��5�k��|�Aϝ3�_t�E[g[��XKA����V�x���ᡇ~fϚi����X�[���q�F��;���c@J?6"2�2Pb�L�/P^ic��:�=mM��8&Jt#�`j�&IL���54ԇ5����}��Z������g���lsSk�B��P�Հ.�+�(��\�RB��0N[��#mR������L��g���&���$
���2 �3�\(�Q{�ya��k��-]��%h��@d��qmQ�z&���-����$��4��z9�j����o���2�8���7�f�݄�6_i�O��ub�GV�*���/��q�5�8t�:�c�����z��I��-�L@���TЎ�*#Y��I\��[�]��� �� ?��;CYY~ع������o���o߾���]qy:jW?>�`���bEbhf&T�W{S��RN���� %��"U�cZzͦ��K͕1 I/��v���!EҔ�t%��}�P��!����O"豸�/=}�\���G'��ZG ��;�>���4U���(w֌�?@�$�5�-;x��~����O�R+,X�r�i�QE�����ן��R�ں�i�{^�)�D�㇯��4ގnϋG��,B�VT����9�燝;�����䓏۹��i�Ĭ�tP��=��J� Y�=q~7�<��o��%�e}����g�r��qM/&�
�R]wW���9s�9s慒��������BWW��������2�'赵����ؾ@o�h7��xz&��'7[�t]����T��&MAq.輢�(wcl����D����� ��8� =u�(��L!�?�r��?((�"~��+ɂ���3��#�Gc��b��Sca�� E�5(��Т��}�p�R2��ڜ%�a�iE*k�?ϭ�L�Mɽ Z܋rޥĈ��y4��� ]V�6@�u�����^Oϣ� ��x�� =;+Xq~
���6n�d9�@�"��{���5C���&k��pR^A�	i`�P�C1X��%NEJ	ԳjLH�������+۳2-p�tͥ)}�M�:���
��q)���h��0��?��;W������}}G����b˖=��y~m%�]]=����@g=R�� $����#�H��?h�;���Z���#��Л�Zl#WL��"	���;�[�󩓝1Ġ���(f��55�<M���2���2ZJJ*�Z�N;=�ٳ+�߻'�߿7�ӖR�=^\R���ɾ�1�:V럽��%d2�*�Un-��=�{yo�"�JOBj�M6Tbͳ���?u��0q�T;?�	�Gjg���w��':����ܽ�`cCs6�;#t�Lhd��ca- 	D�_���<���1���$
 �A,t�(�^$�b�\W~�J||�%�=�L��ǜ�e_�G�QDn�B��O'�)(Y� :���U)N�o�SQ׺O='���������g�cQۜ�ٖi���^*���c=�a�{�L@O�G�/Π��95�"�KMF4?R2AY���z��zvm�Q&�u��1�aH���C�w����Hw�#滿�@����-������JS��ա��X0\�=B�W���|q�m��`�	<�v��6^Z�lT���:h�Q�B�����m���DM�%Aq����iO�0ƾd�X^��"��*H��<ab��]p�g���D�����#@��]���[���������gr�5%0�u��c�Ƒ#�l�҆��[o5�铟��)�P�5���ֵg�x��$��K�gъ�9�,�����J;׋7�M�6Y���ŋ����=^GD�rM�Xp����4>Xc��"$e�%�'�Sv��d� �]�䁌%)�����&���;vXwB��3�
6弌�qY���y��z�d�̝y�
c�P\(��g�������t�Җ��t��n�v����(��n�|�>t	�Ǵ�@��A;BfZ��҂�.K\AAq�{б%"�9�re�J�S�-i�v�ȇ�C��E��96tY�Mui@G�����E�_[
Q�Nz]l�k��i�JYܞ���̝gAZ�k�F{��'��ʴ��Sg�Ė���XK[��R%J�c��R�ilE��{<�]�V|��{��fZ��,�E�����] ��Y�	�(L �%�o,��/8/���̒Q�:�Ebm���Y�rѴ�6����@�b��#���y$���O��xoŬD�����q�nuHY�'�G;� �<UݸV�u�_���o�̉������@SS�rˎ��ֿ������Ck5mifNU0�M"�-+��ը���?y�p������{o�=�x�6p>K�Ġ��^ X��;���_d��x�w4�-0��s/����-��PZn��B������0`e���#VU�R.��c6�Y��qB@�zB�� ��sܖ�qՋx�'®�m�{f����g�
x������9�/�0�3oa8m�PQVj5߉��2e�'������=�UpN	�'�~�`Sc˰L��)>�.囋�~��d|�, ��%kV!@�$	�� ���$D_
Џ'��bI����Z��e}�y�>t�Jg�O�Ё�k�/ڒ.���Xo����2�q&D�*�#���h/@�{�^� P�;�(�"?QsK���7��&]������98���@�RkJL䛕��X����9�8��cʝq�-t�;�r�8�Y�p���Y�`d:�IP����`���l�o��u�c���EϤ��*��E�������nm  Y_d�/��Y�!�9@4q��+/?��q���{��c��Џ'T4�(sP�2kؒ�ʊ��̙3~v���)++)"���w~-#�֖�iˋ{_xqc	.�����{�G����z7�"��ٳf���˿���Ǭk�������Ks>|�gj2��E�s~(w��/~�@x��M�>�AOS�0D{a�w��6ٳ�<�S���ŋ��e�:\c�#�6���}��Rt�?�М�=	�Oz.�F����f�z:���U�Y�h��P���e��q�I�&��BĽ�	���$�ٟ�|9yE����´)S���^SS]�߳���V|��� z����V7�7�'���A �ݭ]���d�Ɩ�nl��i������.��}3�6�-��`���Z��\�q�E��8����4���YɦP$��
��v��|0V=.t��II�RB�E��x��5��{��S�4�zR�<5L �*�)9=]�`��TV��3��L6����b%��w��v�I��L�(^���h�Xaa�Xܪ���~{�/ ��k�yE�ӓ��g�@�"uN��O�})M/S� ���O[�$	VK��dy�rb(�lI�s�␔`�\k�)�eS[�y�����y�<������k���]�k��f�r�X�q�(p���giM�|R�^��JP���FkzV���#7����˗.]z��
�����G��;5����I9�E�e��"(śu��C^�k����}�{_���?l��ȈiӦ������j&e�R��hxV�e=$]1��MS���������}a��-&O���-�l���������
c��k)�ٳ�s�>7�ݷ'�2cz��h3]�9^���|�Ϻ�o>�MC��^�g��~�o�G2/Y�������>z�X���͝k ��/~��/�21j���S�A{�c:�:BiYy��&M��7�<"n�����_����jW�	:Z�����u��[��I[s��� =mE��f�����*��
`%�c0���|���q�U__@/˟�����aбh��ݒ���$RҬ�$m-��>�sr�t�8e9ˊ>�}���'{�
�w^�H%��6���k$��"�����w ��Z�k�^�-f����d_�2���p�e(K[�
���� �'+B��tz�w�/�/M;��e�c�dHy��3$���C��9y��T%�"���\iM��Kpߓ��qVa
��ڣu�NI��WP����tm�u��R<X}��7������b6r�����C�$b%7^W0<���{(�����(ȃ ҹ$^�o�y�Z�t��Z���
���jj�N����잽{.۲y�� ]�e�0߰.ZG�����p�7��~���/)��ϖm;LV��С̭�D���u��`���6��?�z�5"*-/�����i���v�~�Q��������d���/�����֙?>]1G¾V�3~�a#,��]�Xgk�؃�����ɸ��c��K��]��o}�[�\��m���Ǐ5�EÕfgVe�R2m@/*)�-Xhnf)�������u��/?�j��k��7��;Z�,tŉr7�L���δҹ٘��Gy���9���:6�f%e{$�kdN�(uG>M��9���{&���,B���&<'�`~��B*@7a����C'�M�s x�Hhǖ��[t��H���Z�f�%c�s)�YJ�aas68�Z7ڧ�.�Ϣ��:��=��Hi�,_͝�CV&���kי�±�Φ ��8)��Ε��^���H��537��!��ӿ'�N�;s��E��Q�޴���T� �!=?�#�L�:)�oƘ�miiK?3���ɬ�O�w4s�I@3DzF�]�^�o�i� +
kJ�Xy��J��A�t��H��0Q�Tx��Q#F�bg���{�YW�X�bӫ@'��͍���[�)**�K��7Zp��mj�T�(Oe���b�"Ms�S#��7{�,�v7m�f��� ͭ�у�`�����$K��K>;�tƴ��NP.���n�M���%��ӓT������:$�Yp�Uׅ{���a��m�&7��Vkd��h�eX�ua=�J�Ñ#��~zY�I}��b���Ś��r�)��sӤ��bx����0a�x��t�Cf*�DgIiqhk�ٹH!�?1���v^J4<8fܨ������^�
yM��i˦9\wE&���9���+ ]$��}�Q�3�6�4	:	G��5r�$�.�	0%tcp�y9'�b�g~��<E	�E��w�i����R�;��F�z1�k<b0��H����#�.JXZa<�:�1B#�b������ :Ѭ��t%�FB�X1���O}�9��v�8���8*v�B���P���x��wdX��R4��^|?1����:�e��EK�W9�n�S�>�C�{zV>�ŁE�0��&PA�*&�a�K���+ `u��}}���!��qm��\�N�{�Рh����}��W����
�͇>lذ�g����e˖�{5��䱿� �yӶ][��ǳ�֭�֯_oeHP���}�]Q��&}-;茷�
�N]0�������bƺ�%F��E�x�a�ry�|�䥡� .?ש�������	sf���Y�.�#Z��w�u�L�_��K.�̺��ڶ��>�q��+�1lXE3f\ڢG�nN"�9Fq<��^w��H)����=e)z��8���F��n�-���?m{�����'c�9��j4L����RK}��`�;Z[Bmݡ���k_^�jV�k�-[��s�Б�_�BW��KY�>:�/�O1zt��R��l�P��Q�� =Ӈ�R�.A,�(�fq�����v��S)�\�,J�*eMz�~<@g��)�D��ӂ�p�3�)�lc����x*-)y^/�@?oƩ��!����E܀�ĉ�-�E�-�i׈j��1hfZ�R*������9/�u�x��3��/�`FQ�X���Ҕ3�.�D��u��osp/1�:>t�����!�]#��Ȼ;;�l�@֩y���M�����Gi�ꍂm/���,�f&)������8��\)���Y�+E?CU���T���6����& �4e�G
hQ>����-�y9l���~�{/^��j��c�#�}Ͼ��|��o0��0!lݺ=<�쳁�z�Q~����;V,�w q�(�k����@��� :inX�V���Q�e�����uOa����K��`�5sv�ͥLGh�1H2v t��.�L]z��<��n>�9�{ �2��eč��&O��r����8<v��1ÇW�w���A��>�G�{m�
Ǹ�jY^b���kX�Ծ��?����}�X�_��?�SW\Vji�Vsr0+̘1+̝;/�3�R�h4�7]qƭ7]�������;v�����AK&�n��G
�Vbl��{�[�w�!�E�
�Pp=�-V>b��$��1�>�u���.�N���qԣ&�@)���Z�t����y��؇n�X[�ip\�g�5�[���5m�$?�rb@������� �KB��J�+�4��7�7�[�DՎ=�";��BcY I�B|��Y�*%�@"Z�����X��(XP��?��Yh�h�ԡ����I��5�kd�z-&)h��t���~�-����q=~ojl0�Zc3ca�,F�G��&��x� ������q!jؾ�t����J��p_z^X�J5t]K�;�ڃ6�ɺ�^�}���P�祌9��aÆ�6b�_]{�U�}����q��x�߭������=̝??�ڵ'<��㡲r��NooO����@�%�:ۼ�
J4���ed���,��]�e����85���4ga��9�1F�����JY�l�a����֤��-���!P�X��\s]��O������n���U2�=C ���6{�'���RW����:�'<���L�2Ũ/�1��t֡���:0ФgR���_X�
z:�(���3�Xs��!E0�o�oЛ�g[�xI�1c��GsK}��M}�������ҕ� }o���V��g��>0�l���VP�+����׮]k���@I�Ȅ�Z�%�NeY��s��e�c�UV0��ye�e����j�c�+� ��cʝ4(w�	@)Ct���b�<��T�Kʈ�R ���ig��]�6�C�ORBҚlN�m<��L0VB�r>�Ga*z�@c&�ge�߲�9wo���P��*�H(̡����L"p����H&�j�����>��7�d�P� �k�C���/�K���^��������4��2��k����&)b7x�rqe��[G���lU�U��X +A�C�e�}H�E�f@���u���wyvY���\�E�
�`���Mi���4�=�S�������o|����q��H�RO=�nk���ӛ���Yg���
k֬	��^�D)_2n�C0~��b���9�n����{A��R5k?t�*}�:���e,c_P�B�|
a��i���<����փ��nJ�%{	9���iӆ����.k\WE���_hSʳ�ù���/}�7jV�뎿۾}�KKʋy� �yfB��p�	v��#�	V3%�ߔ��\S|�{^�"/`���1I��(�(3꽷+'̙37̟?�b�:;[Cu�����������	Ы��/ݷ��g zk�kx���]�:�*����G-�b��v���y�,T��]�K�
�M@'Ĳ��W�-�Y�.  /�hw�/�W�s0u?zOW�-F�O�&BT>Yʲ�%�%�m��9Ejc��~�8���x�1�o6���e�8�(�O�S��y���gZ#\"0)�=ĺ���';��X�*������x�^pY�E(����>lxe(*,����z���y��GL!R9U4ϣ��C�ruR���^��"�p(DƕI9y���>��wZ[�F}L��B�g��eQ[M�<�����n�e(�sJ�-�TP+\����j�����J,]s�:P|G~����畿恾�#*�%Q���cƎ�Ҵys�}���*���e'���յ��u��-۶��p/ӛ�/��ǟ]�$q@�d����ZNuCm��4�w�V2�u��=��Л�[�z���Pt}�y�2u7�)}=ݶ� D7���Y�����.s��!���`X�\�2T���͛6���}��W���T�Lc!eD��q���՟��i�2    IDAT�.���vs�5k������_}�hu���Q�6n�j5�>�z �<�=w���aI�n��]���x��_��s��EqOȼ�P\Bυ�@u��/==�9�hw���|����z�/_�j~M�^SS�h��}������<��k��4�n́��S��|%%\�)�lTV�@]Խ���Y���I�P��⎹6�EFP'�d�I!H�b�DZH��8�\ik4/����������n������1�p< �)lq����+@$�N���f���I��4S��(߬,�ȯ���p�����}{���/d�!�Θ�[�Fd��P�t�r�r��aWgG��h�@\,\�������lp�[:���;���;<X�X\X�ѱ�-�ß�;V=��D��4�%�t	�m,�h�5f��E��(�(�)ʖ����՝ԝN���>�e��R&ET�$�$Vp�`�*��{#Z]tz�6����(A~G��(^32����(L����$8�qh�1zԨmcǎ�܌3�9iҤ��+��o�c�����C��~���n��&+��u�{\8R{4��]�f=��a��v���!��Ǐ�z����զd�^���$���a����PC�h3����6b�Y���JIY�+�!=iw�d��Y)�_x�ᢋ.����h�|�?>���R�y�6{��RÂ��;/��$/����'L�6�?~���j�����ԯ��݇�,Y2��$��/���{�zã��	��u!+E��� w�D�	��s_�ɎE���}�ږ��Wv����QcF[�wK��Yz�ƀpڐ���{�����,���uuu���~������Iq/d����,$ =Ӛ6p�tL���V(�7n~��t� I(���#A�<kY�
��=�ߓ�H�����gPe��g �ҶD�g�zNAD���
̙���.�tY�ڢF�g��% �ye]�A��wc�Oʉ�)9:&�`eճQ�:����o{˛CA~n���1J	�7m8�-n ��UH��b)s�ϳNI�gM�@>�J*�����} .(:�l^9��6�e��1���� ��aÆ��SO�`aL��0�]ݞS����z��!�>�?Z�.ǚ���"�P|T�z���$5	�L�0<C�Gs�u�I��hP,"gF�������m��ֳUo������ՙ��wf�
iRT���(�{���M��w7m7���M�$��Ĩ�D�{�7P:(���2��������r��	d���}��53�~��{��{��y��y��~�z���(?̹�~-G���\Vfz���w��,-++��i�NJJ�-��^�3����S��b
�45���ݕ�ݚ5kܦ�[lm��Z $�y�I3�۶-��@]���>���5�4�ݻ*l��n#�
� �?\�&S���*/�� �u'@g1��.k��&��?gΜ�ysfL.))����/��'�l�����;v�u_��p��[O�OR%D����2����6�p����t�M���^w�u�~�g4�|����Kݓ�6�e�i�����f��/+��-��%�^���5�x7��y�k��m.3;Ǖ�zbQ����=��mK����O9���zeee�����546桙�ҝ)��5��{|�8'@Z�!����D�)"`���5.]9�a�;��]1p;GPu����e�`��!����Hq�/s�/��g(�V�D�:���]�.���q�_�S�.�]��<�L�4�R������!�� �����X��eg�6Ӭ���2�4���ޓk�}������`q�*?׾�	8�)
Xs���,�d9>��b�ca�8�4G����\��ma��.�k\^,�����]]C�#nF���R� c@���/���q,1D�������`A��2zh��6�Ĥ8 �Js)g��sr�\S	(��о����"&�'?��Ph���e��	O��5큜�L8f�9b�(d���7`���ǏǨQ����n=��̲Uk�ܻ�zy߭m���sϵ�'���kKm}P�*kv�R/������[�-�����U�ָ�}ծq����j���sy��]qp,t�zv�*mY�v]�*���~���l�_,�<3�j�Ϟ={׬SO?hРV���֊U+o�ڷ��t��6��gX�����S]a~�knnt��r�Y�t�<=���G�����o޴mr�}W^e{u����/tͭ-&ۖ,Yf /@7#�B���ǐm���u=F�n=��o�0E�y�PdJ�X>�ef��~mm�0ņ�����U���M���w��j�� ��/~��=u��N�&�J�Z��� N���Ԅ���x�?1���0ެ�C���p��q�,1�̔�H@��H���)��h��BP�<.^	R��*��lo5�1/	��e�'��C���C	{����З�EZ�!����}3.q	,��ݻ������q'�t����<p߂�/����EU@�4/�P8h�+*,v����	'Y7��˗ۜ��c���r'���i���  ���Ys\aq����+H\�����z�rح^<\�u�]jT{�����p-ں� ]����<h���dY�y}?Z��_���Bp�}�7t�"X�|7#�!���M�u��-4���� �D�aQ�=Z�0��j�LOs�d�:t��ƍ{�������F��?3��Җ�xcG���A(�m�-nƌ.7?��ŋ^�uþ`?йC��7V�1wvg[�zQa���[i�S��mU�V�(��0�ꪽ�p�(@.�9�� @˳%#�5���f�0k��W^~�ؤ�$��w����{zwE���;w�{M�����6�y��P��wv��Y�f^�?�WO��W��K�W�y�=��b{�u�-rs�a��O<e��^�����BVa�Xzo��!Mn���X�|�^^��LrtE%e&ךZZ�y��@�ќi_U��5c��7}���i��ŀ�t���յ��e��0�#��X�H�����1oɂ9��	�aU��S�dY�!���:͏��B���t���<)���SnlY���B
)�񉭍�����7t��>�qO�	mƠZ�t����5V���H�u�>v�<H!2��<�C����c9�,M+���@r��Qn���f-rL^^���7�]g�g��YRRd�Tl���ƚ`1+>znJ;����Ƃ���>`�c5�0\{�XZb�\��f#A�Y��k͝^�(�������1w�C��׻����=���7ε�5���l��=+(��\"��1�k�z�:�	��N����ƍ�MʺC���A�(��+77�#/7��1cF}gҤI�H0�������k��\�e����,<��1c�s�ƌ2��{v</O����<9��nú�8]�m������jn�= tַX��)��)�y���2@��mi�1o�q����E��*�\�,f�Ҍ4o�ϙ��K/�ĉ��k�-?���^{�����.�쁊��
�(~�_���xF������-[6G������я<���{���J��6 :d�y6^Y�؝v�i&W��c�{Y���ȥ�
�<��׾iq���+ג�-�N诨��<��=Q|!���@��Em]�6h����߸�V�_�k־�@E���+��fd���~n�� =�.<�-[�Xi`'N�E������.���V��V�YϬ��x�:O�&��*^;�,㰰Lz���U.}����θ{@�8��&Z硕'r�@;QAJ�������PQ�s�\�_�J�&�3�L���!��<=�SܠA���;Zi6�d�kӺr����v/�O�9��y�rs��&N�d���qz d⁌˄�U��+?�d�y`���ifbe�O�R�W�z�c�l�b$��2���x4_���&�×����#���Gy�(��g��f��V1��B�2Iq
�!C��^�w�?���6 9���_�i��Ҳ�ߍ>��c���N����ػ�v��;߬�?`a*d#��)3Nq��lt�-^b��h+����q��W	Պ�{��X����[����T7m�4[�b���v��d�Α4g��(��wk�qނ�b�݌���s�;zD,�7������cO,���o!몦���Ϯ={\����n��p���
�Y���N����v��w��ܺj���445�ށ�@��E6��jmm���uJW�x�f~ #�>���暫ݲ%K=q�%Y���C��\#��㏟8�w���2�Cvj�3w���xh�p��/��[7߼}�oQ�!
�-�yKI:8�]�*� ��>n�C�e�$��dፄ֥,����0��;`߉�z���ƽ����j��f�1
��"	Kil��C7+��˴=��6t�m���J�����5f��Ρy��'�ax��%seG�n�)22,�̋�^@���C���X\�` �w6n��:{zmc���32�sdIsm����LOw�ƍ��p���۳B@dFMcZZ�}:X�'��#��sϻů�n�i͝Qڃ���
-�Н�5��B��|��Ø�~ld��q!��e!O��>��+��� �~��{c��+4����~���Z������Ҷ���E��(֭�F�z��������F�3��r�9;w�y����mٲ� ��5�yf4-_������!��Dd��o��[��-�N�n��:�+� ��
�1t������]�.����j煌����^Tb�\)��?���Nv.�Yk�w�y'$��ڵk�_[��Ɇ�ƹ���:���j:���\"�HsK!�BH��5+���n��+3���WP8������ԩ��kX�Po$��_��5y��d�6���0�����^x�9���r��������[Q�n�p)�CM�54z�Иqc��Aiimr]mko��'N�:u����X1��سg�֭[���'���� �'�Eݨ"�(P�n�M��;���E&��Z�c.�.:/��.wYi�������L���tΧ��YP���rL"�]ָ~�r����RPH���>� _B^ ���w8�!�'�g�2�s�����! ��]�>��n���ٔxV.��|�aQc���fվJ�T9'u�鲴m�s��N���B(/Z.�W Z+�گ^�kKD����]�ȯ�|l�k����������֑�ጮn_�%|IӖGB3�!��Y)�Q�Ks�u�=��D9e�p�Ӛ =9*0!��t�!s
�ct��*c�zNf�?n��=��G���͝{��A��3�;�?���G
}��ߙ�={k�ߵk��-�>�1 t��X�����Mi,2�d(�ì:r21c �v���zb����f������d
j�O{������4��@y89���Ξ�;��E!/d��B?k֬�����zR���8s��Տ8p �x@!*�5�Q87��~?����\~���~�K��4�\�`A�=�޷tݺ�̲O�\�md���d���/�sZ�RRl~�ir��w+c���������_2E�3���ճ���r���C�<�v��Q��36?����@S�>��ɧ�rJ�ۭο�+�+�nX�yڅ�e�}P�[-�e����⑅k��w�`ɒ%��e�n�VR������ka�W�J����N�otm	o���;"�������J�H�j��a�Q��-Q�:0Pu��A2f���6��RZ����4F�}9��y~�4�qEP�$�-��D��p�`cN�u�O�r������q�����KO!��c�n<���r_�2�zćժ�j��k����uTV��h
�}���(����3�O8�Ds1>���V�#�� ]��5w�KݻY��UkL����d���wᅫ�uH�]���4�7}P�����Le�i�#X#����(���<C���Ӧ��__li{���]KN<�ğΛ7����� ��]}wr�زcϿ���X�Y�xo��=��{˦�B�b�ÁX�� '�GFF��2�`�k�듗�e�&!E�G\�5[�5��F�1�H|�����b{_t�c�`���伨u5�$+],wR��̚��%�?�pO�7z����2���K��c�V:�V�?߼YT�����嗞������~�3O?�ܭ>s��Σ4�~����w�u5�&E��!��&�+^fed��>t�ۺy�9|��Z�v��^������J����v��c����564t\õ']0o��c
�.V������6����F]��|�w�HY!��-PA@�(�]�ܚ�t�)�pP�{
<1L��kC��j��X>�J18��]1t���R@�.wz��U錍��D��[�@s.݃wy�0��iY�K]�:c��8�c(�0{��kҼ�6;U�p�g�Qk���N��g����m��Q+������ƯY��Te�B�;�Ć*.,4AAQ~�|�xR�(v���wܶ;�.�MK�4łz��^�FC�g��w^ܧ��
�=���1XX2K����=D�(@o��NW/��u�Ÿ1c����) �n���͍�M���*�7�=����ǯ<�R�}0�{�n��ݖ�Λv�4��}�5ܼ:�V,�4O����=�\��w��Ǻ������|A�d_���T�Z�P �J[��NV� �s*���t�]�k�BGy�5k֫��?��=�e�V��q떗�Z�%�X�������G�⊊����ֿ�v��g�缿��/����߾�s��4J+��>�ˠ/~�fSj��l�*�_A�1j��M�y���о��u��GܔNp���^))�Q�}����o �x"�� z}M���+���K���z,K_�t��U5%�(1+&}1V�=����D��Z��,9����%��nDBVqiq"��X~K�T� ]� ����x�#�����5��,}���]�AYS-|�������5Ѧ������F��ɩm��Fr��CpW�6��� O #�^������2���Lo�JD�X�J�˲V��kaߍ�Z
���\�`���N�@>�9��4e�	Y�\�9C 0'�Y�s��,v��gq�C��{��D�vcƌt��mr������W���ɡ���8T,���f�L5ϡ2�P�\������rm6)��w�<x>�3�f<X�mm������7|�0y�Dsߙ֟�s�G7����y�s�5d��߆���{73�i����7}�@c3qb�g�oA���i ����^���~����lX��*䉌���b@�����9�.�I�r�o����{�+����W!ű��K��	͒a��t���SO]t��g�|��X������#����{ｮ��.
�&��v_x�=9��̭[�֝~�iW}����[λ`���G}��K�,��2�܇,�~�#��lڸ��y�yo.\��v��T�Ls�y�\IQ�N��J��/��fL�ic�鎗3���"������c�wt��_x�E��p���<���ɗ�\���b�x_����G)k��B�$�-r_9����}��#����{�I�+Ʃϴ@d��!��� M��R4k8��s�}�D��Cس�DU�U`�uR�-�� W\n|G`�{����s8]�*�%Б�eZg�A����Cp��ߋ��Ey8�w
)�7���=#}֬Y�[��La{G���s �0�ॢ3ln4c��qsY���d�$�gs�̱�z����M[l�!��7 �� ��<J������ӀW1t��ʎ֣ kķO�����9�5箚���3"V�\i.R���#L[y(�_���c��ޜ9���/���������Y��ֽ�5�im�0@oh�]�vWV�뮻�-~�eմ�z�@G�hj���J&�nW�\a뒸3�1�9k�'r�Tcs��)���s��H�Д��a��FVx �/��7�$��+���&O�L�ܒ�_z��VO[�z�E�����4����n��->ݸ�W-,�������46>����M[��_�~ٓO>�pu,\R<dw�E������USPhF���m�.ʇ6<���nM�������b���nr�{�[�q��$0�;�KIG ��qD��u��sξ���_�c�׭~t�ΊN��y�r�c�3P�0�    IDAT�K	c�, n��Q��tr��>��]�Ԯ�~�\��e��A����0��"��B)N��l�MNy��CP�1�nt@�Z�<8�o'���"�	hCw��F.z���<t��;|N:�ί߄̕u
�ZƼ�EV7a�K.���廴4*���piyw��ϿhLX?�>T?\�s���<�|�`c��o�.���	H:|�M����gźl��<xb}���s�a�»�}H`�[������+q]���|!$T�B�{�:��̰s���q�w/xЎ��Y���u����.8���s�ر�^p߫o�f�����ʪ��$�`�Q��ZW�o�;�sܦ묬kMm����>4��>�'n
3�o�)���V�}�P��n@���Iѝ�����b�I1ۧ��M�D�9�!@WaR�Cǳ0y��W���C����x��E�MM'��g�_���n��K�u$8�}�le����+/����5+����~��~��roU*�� \���|��&^y�EtC��9��-�<�X闛�9����U���}ν�����+�X�*��\�ȐoX�@�ݦ�����.��������훿�u�Ѭ���6vQ�y���q�{�=�f!G�y� a������v���B@W]nY~�>	����{t�p쎳��V}"�3��=,,��r����j*�漜�1���,��j>�����*��������ϲ�oQ�|Z
Us+��ax�#ז2�F|��WFu<(�e ��r�o��d
��2e����NSk���kpy��LF	�sۍ7�h���;�4f\�/�H��wvv�)}�;�+)jz�X� �㒕����),��8�2p�q>���<ĳ R<�a����s����]�~�.� ύ>�ћ���wO�0�>�[~��شu�������wE�S<ٴ�j�[�j�KO��A�KI�5H#��!I��@�:��:i_�WVVb�z�>ߋ܈_Ç�K������Z�(�(X��!F�*0(��U�X�Tv$�7~��eW���i�4��m�pm]�T��>��g��l�$�!@��N�ʅO=Y���}zڕW^i��,X���?<���%���{��8��_�j�3^x�Y���e�1����F;�����G�a<���3���;w�yn��M6Ϡ6�10LR��\J�/�ǁy#��|�ѝw�9|ຫ?怾�r�u7l��J:�v��G��<t�b��'H�&�a�!j`�Ȓ9�%
_n�&��xBw|T^�{�<nY����#őz M��k���rOtb��@�[�s����<�ZrI�;t���r���9�{06�'	��@��.�>�bވ��^m�zߚF���l^U:�|�t�	��uÆ��(2�3܊�,�P�Pq���5��8�nT��c���j�̞e� Y�0��N�Z�y>��r��-���� �wg��V6/�f_����(,"O�s��I����ݗ��U��~fF�mڹ�}��G}�]zZJwaa�3g�����?����$�{�������[+�klj:���uL�䪚��#���d)e��$�r�$eI}a0����i�F����~P+�B��(-��	�q.��t,t��	�^6зe�%c�1p ���ѣ�\��KޱaIuuu޾}5˻cn��O�����ȏ*(�fg�'���\��M8���o���2�_��o��?}`޴e��7o��5��p�B�l��4�6�d��u�jBc�p�D̹뮾ҝ>�4�����H��IO�4@'מ��� m����]|�Es�����9��ڻk��-;�������Ԗ�%�{TX&�!)� �1J�ܲe�L�3bYd������&��Y�"���_e��(C72Cښ4)�P��Z�XF�-t��[�@�Oٹo)8#��@���=N��%@��˹�\�6ƨ̬�]:�׈}�]�&��"v��E�PHB�����H$���TC��<�f��1�힓SLk�rX,jH)y�r��٧���>����uI�έߴ٭^�ҵwu�I�Op{�W�]�w���|7j�����R\��ܷ�Z�9�HI�wkK�w��^���Y�h���6�B��9�`)�0����E!󆅎b���z9Qk/��Lu�>l�հ��L���p�5l� c۾�꫕9�9{���9}��[�Ν��]��C�f�����ۖuv���/���%^�-�����&���a lFV��_�Y�Y�c�\2� ��{zԽ��Y�������r���ejVz��S��7zi��*���}��r�)��wkx��n�̣F�Z|���8�G�e��ڻ�~����'��}�،�گ������qc]Kc�������w���:��}�_~��M���/W]u�����sϙl`\x�s�}m
������7c��,�8���w�\7}�4k?�A��n�cSS,�9����:]9����']z����9�7��׼�fGm}]�
���p���֮k�8b&+��
���"	dD@������4d�v:}�>]')��T��"��f��q�a�c��2��@�w�������-��4�x��+���o��g:��-�/w�<!���P��,eA
�\\�GC����c�ÑH����]���k�3��͋��8!��s޹�N����6ltϿ���<�8y�+)*��ǹ�9�a�[;��|���<I'͊O@z��(ʧ�:�>e\�>\���WQL��3��p��87^�%/o�G�����,dވ�v����'%h¸�& 9���Ĵo\��^rѷKKK�jmm�߿��>�����c�ib�X��m�6�uty衇�����d�.�>@r�X�"��>�{ ;�;r	�tYü�~�b�zGn�s��-��{+|��N���n��wˇuy����!���9�5�r��̙3]iY����x��������A��͏��[N\�~��������R�>�Q�*-5�Hh�I�T����'����;>�������{��f��x�����[�+�LS����8�?��,����	�&����S�O�9��8Z���g8�.�����͘�~��ڍSS\X���K/}�g�m�����L$�R�,Y����zxK�Ǩ�uG�?<n��.+P�I��������o�����\O�Z��kO��Z�� �� ;�@=`��$ R�9�I�^o��@&:�YqR�MO�:$�SB�`���=������M�|�טu��V��Х�ȫ!�NT|B�>�޼$Q�\��Vz��v���Q���;�̱���s�Nl4��5�ML����:7E�Фt���n�ѵ�j�hc��A��v��qM��	Х`���������)�������F�8�nv�����v��S�i	O��p���o���b��u�7W��H���g�龪���z�$L5e�I��-����ecr�屷̵��g�)<��q[gG���5 "�R�Y�tMd�pm
�x���Ғz]Ww�+���JJ]vV����ͧc�zy���fg����J���_s�YG2'�X,e��Uw|��_�YXȵ��FWп���]��Dδ57�Ԕ������?��]W�����]�~��G��O�.uȄǍ6e��ϽA=��y9�>t�����֪�~��k(B��%%�������e�2���f��N
Lչ�%��?��kƞt�Iow�Gй��ի�޻w�Y����Q޶ =n!�S���3��b�6l�I�Jt��C.P
������L5)�~"��|��4 �<'-b����}]?�z��G�B��\[�� *�ei�y�Z�rP�*-f�tp������ga�A�\��I���(]�g-o�&i��LT� ^�Ș3�?J������)��F.yD��z�gC*H�o��� e΍�����oy(�yD	�[�A!Z9��Ç��0�1{�af.G*C�q�>w�=���egg�3> ���������'cƌ�s��эG"���雁w;{�T�����]��-[�&PP��ď?~\�[�?�)�_(�V����r)��E"�`&�����r(�-��
��%���;�lgߢ�Tx
 ���W�b]�\�ݾ�PqQ��o��hĉ"�F��0�U��t��>�*+{↫�8�H�$�%�����K/��d�Z!��Xt���%ǜ�<i��h5c���Ӆ:�m?������~��'2�S�]m�g�gdg����c��{��Ǜ���\�?�RNǍm���O}�����}f�wƺ\z�^���M6���Rռ Ԥh9��._��������;j��q�Ư��8��y�, ŝ���v����]�,�8!#%��ܹ��A~�b�6e'Z�:��3���@' ӹ�`�`8�&�:���P�nĵ_�#�r���`���.Ѕ�X��d��@�k�>��NԦOV����E�����(,!�Ң��إ iN�u�Z̅����〞�����t�yG�j����A�� �JgQ�ڬ���q�{��R  ��xg=�z���+qg�P���(�^p���V����#�5��/p��Zn/�f��n�ر���d���þ7v��Gt0�x$R�x3P[[;���j��-��E��Ϋ����g�p�$w˷��$�e�3��3��}!�VfV�������� ׼)�j��#���3Z|ȫ�mߺ���V���2c���.2� �{W��f�%%�����^w$S�����'?��� �E�^OO�����nt����:��|ᅧ�ӹ�,Y5�۷|�����A�C�^FfN��ã�w���lU��)h�u O��W^�.��B�s�������m9�=�I.7��0�d�P����qc�����|�;��Q��;w��m۶�i�'@P����_�V�i*K�!�
��D$c�q��p�D@Wsh���.kݻ�}z� [� 1��BOT* �	Э�L�r;=t�GqpY��1,�.P
��t�����4n͙����6���E���]͟���c���2]��$��ÿ97��9�.�N]�{H@�	�ϙ�*�� V/�Z��UO�LIQ����O��L�0�9$��$GIa�2Y�e���&N��Ŕ�<x��iӦ>u��S�����g�;mȾ��f�h��ox𱧞���۷�=��N�9�}��u{vWZ�T ������V�#�sޓ���tMuܰ��(���V%-�a͘R��8�e�� ��%���6	I��~��fЬ[����l�Ⱦ����<�����������W\z�?��\=��3��z����b��QH��p�-E��|��l@I��ڷ`��{�2����O��-��j��'�(s]ݽ������G�p�c��؃Y[Ə5��9�C� ����4��4�fi��Lq�����Vc��B iΝ�����������~�����^�~��ꚺ$:	i!��, L��`��L8m��L�`%)���,���]�v�C;w����tҗ "N��!+T�.�� ],} ݀ʊ��ĭmj��b#��/��F`.e TjB�\��؉����Y�s���4=#ͻbf���S�p`�1�Ѳ!z{ͥ�K������E �$j>lQ�kX�#��<pͣ\�lh<,X($���s^)r%�v�h��P ,{rWEz4�&٧Ԝ:�˅����2dȮ����g�y��z�+�i#�}�7Gk�y��+~��?��j T�<q\͗]v��ꚫ��T_w�RC�M�=�����Mx+��_�1���N���;�&{��ʾ�諎k���#w; 'Ä�S��9�Y.3+��������0Y�5Q��t��P=��3]QQ�/^v����vs��#OM�㧷�WYY9��:��gf�˝X5)c�d_7��wm��Ξ7o�uW_q�O~v������I���"��������R������$d2��������n��3��/��{��=�?��rsP],��4�����׵�4Y5���;�����Q�����ݻw��_S���V�3��-�9"���.ДU% @���u{e��;a7�ڥ8�:�ib,X�fDqk2�y8���]@ z���̧�%����Oˌz�B�ЂH^!�'�uh�4u�8���Ү�Rb�8qκf8ϼ��s�r�I�y�b�Ęy��e�=��°K��M�b�⹮�Ii���U� ����VT� � t���D�&�nyf��N�����nk��9�X#Gx@�r����g�uV̀�������"++����т�����ڵk������7l�8˷�%[��~�]r�%���[�.q�͛6��s�z�Gl��x���f��* �B�y�V_�����Wuuv>�5P�ٟ�T��{�/Pù87Jr����-z�G�=���i5%d��n���\Vv�+)*t���w�����������߽�C=��7ZZZ�W���N 7r�1���Q��}����������\j�SsE�2a�	f�ﯩ�Է��v?�|�A�@i�9i��D��~�Yg�&LQ���,��ـ���B�1#��Í1t�G?pݔ#��5@gb�/_�~_U�8Y�<���,���e�CSR��ڝ���,KK�$kT����Dr^�,td���ݻG�J
;��]��V�(�l�3�ut��)~$��� �Jeh�h�r��e5
����r��XY��_Ii��,`�J�;\1) ��9�J�rl�oY��7$�i<r��(qrո/6��ӱ��z$�lՙ-�
h��ƌ�/��yݾu�	-�HL���MFfЙK ���Ik�p�?���!8�F�NJy�GH,�F����;�cIII�G*x��뛁c1��ޏ~�ҋ/|������:~�s�5/`C}cdY6XI�ʊݶ�O��n��v�i�"~m	iJ���Cb��fh�,����7�����	d��US<)Wa5eq�q�r|kV�1�1+'���qxz�(��wFf��W��?b��\x�=�s���?:g�����~��9j��=PoD�,yIC��*�9�|��L'7��s^b˧ONu&M�R���)Y�Ϗ/���q��ڤ�ng�x]sՕ�?����W������ɱ�s�����t�̴T+(����&N8��_����H��Q�իW?����2�J��r��,���)�E�ZIΔ4GqZ�	hB�V'����= ��ؤfpTTF�	]�X��\}7��Éel����yRSlA��1!�������}b=�[�g��Z��<�`������X�|C����9�� +�P@�f3m6*0����2��w8��hn5�Ђ�]`���s5���v׮]k_g������{�7�'�̼�EBq�F`eeg�K]�<,`�3�|�������r����ѣ�
Ax�A)��K�&M��	&<{$��8�3�򵕣���[�}�����4z�x�կ~յwtٞ�ܦ�6�f�
�{��3f�pO<�U9��q�iNf������V��7R��5 {�}��Ki�����BT�Mơ�Ţ�����p�#�V�g����p�Ʊ��Ν�ʇ�ؼ93�����?�{��G�u˖-�S3�3%۬I{�)&�W��nA����w�vٵ��d1�Sc���&皛��@z�-p���q�[�y�?�8�`�0q�y0P@���ݻ�+��U�:���c
�0G��C�7��ƦWR��͞}�̫�wɢ#Y;Gзn���;w_9���~k/�ި0��UV��kY�hD$���Ů���<��zK[�[ ]�脤1�~�.����*C���Ԕx���C�{R�w��]豞8�����ޤ�p��3�y?$�)���;@�:s�5u�<�,Z4א���GaӦ��*w��z؉^�P��=��^~�eۘ -.�D@�V�����T4j�csR���RV����菌�l��ʋ/��Pjl�aÆ�0�١C�~ʔ)�d����d���7Gy������ɧ������gͷ5��SgZ\\ޫ7�ceW�]۶�A�Z�|���aUN�t�ϭn����j����q�[Ռ4\�Ş��FyV�& ]���D^�]���e J�$�0;�����O�ǯZ���:��iM�ͯ�?��<���K^_2���mbVnN:c�lz�Eu    IDATs�=�ح�|�5��-��}~?I�������j�O^���s��� `��WS��Q�U������t���u��Y4����я~���O2��˳`,-m���P�H����Ȭ;v̚K�?�ԩS�QV�Q���ʩ7mYʂ��N������<0^!��)�� @��9�e�	�rW.� ���QA�,:)�ti�!)Nʈ��>w�>�)q@���jIX��N�5�F��NL�����Y�ع���Y�:��R|�@���J��#��R$R��es�l�V�dl"6��	a��]�����b��2N��>��ZdS����fnCoCh��J�̼���xN;`-+_)p,�Q�FX䮻�r%���0e�С�&O�|/��&L�w�eq���f�/��U�6��+7/۱k� d�ǐ�Y9�Ҧ���_�&L�dr����^�t#�m�{��<h�P�#�	/#<����+v�v+W.w�9���f����d��-b����(�%�e&�a���gKr�}���N\�x*I>]�11��L7{�l�����\�s,d�8�~�`r/Fh��bd!������
����x�I\
|���6\�\���ݧ��G�Ƌ�n5����醖��(+���.IS�_���9�^����n���N�,y>����VWRZ�N>a�|���֑.��
���\�~g}}}���j�_��IN +�,5�.�ISm��3���E#k-�q���!�K���9�B�@7ЋB:�q��v�W6��x(@7"D�g�ǭ�dg�� ] ���s(@�����n���e/�x�E��5_*�*�>TV�%`��C��14L6��<2�ȥ81����k�^m�p���/� V9
�96��6��QYs�El��.�5[\.+�-_�,N�#���q*\hy�YF�����RTTT��ݹz�ĉ�L�2�w��t���︾8�3p�m?����y��&wSRR���J�Sg=�]t�%�}ڸq�kh�s�++�}�����Z�*�9yL2�:;}�Ն�������zzq�׹��^ه�FA���\,-`�!>.��MF@ )�P������n��W�MWǸPuP��.ri����׹'d���'<\-�A��7$7<\�|�bojj�G�����G�de��~�; E@g�����_���'�8Hss���#F����f�]��b�5��?s��ٳw�z9���EW�\����j<�n�.o�]�<,	e&E�jp#X}�����BK>%�;&t��e���k�B�X�:7��Q����,wsۚ��7��客2���B3�L t,t���+>jØ�c���%.�G��*����5_R��.���s���v����8BD�6�+%�P������6Z�W�����Мъ�����a|��L���BW�Xa�1?7�\h�+�J�-�ӧ��]^^�f�֭���ӟ���Z:{���G����뛁����G>��ʕ+ϡF9��@s������|j����!��\`�5,붦F�u�3��WC�y�9.`����+��@����%K^w�;�~�H��O�ό�ސG���o�r�+��������n;��*�q�������=��۽{��[H=cl` �����f�F�v�Lc<f�G<%��}�O!f�Z���5E N�E�c����2܃��,�MU{������xn�<���.B�HOf��i���f�h��(/���o��M�fMu@ߴi�Ov���I
�����@).U��KiJ,Jn� �y��]��KG ��,��H�HqF��S�,����G<�J���>���[���e��R?�8!� ���V�\ ��p��_��)�L�[�7�ǅͽ��}ڳ�RMT{��x�9cQ�K?����& t9�ڈ�.��m#��#*h:�g�\�e�BGf��}O �/�vB�&>�/�gi0t �@k�a���egC�?=��=|�W�ϟ�����mIII>��ꛁ��ؾ}{��>��5������=ppyΏ�S��y�坳�7n\�j�ݞ�ݮ��ټn�O�Uel5r}đm�m���%Kv�ֿ�ּ�ܚ���s�Uu����o E��5k�r��I!��b����[Yfv�e:QyR\Tb �~��7����5ʷ�f�#�Pj�T����1�E���!f>eʉ��f���y���g
��< ����=j�������y!�+��d$-DQPh�����~2E�R\y��]g�?�����V�n��Q􊊪y6�_�dX��C z���C�
��Q
x(L$S1c&�P�(��Q
B@��-���\�*,#p�W� =T;��"LI���C@'�.=?'��3�i�Rc]Anl]S���!���4/�Gs&�($��8���_v�K
�@֯���[6$t.�#����a?qa��N�KP�\�P��8'����ϴI��ͫ�8_�"۪������|�>,��[zZJ�ȑ�z���}Ȑ!m�f���73���Ϗ���yESSSVW��~�UWk}P�`�o۶�,؂�Bw�g�Gq˖M�n��ڿ���֚�|ʌ�����Xn�!#�#�?5�hS�Rݾ�=n��W]U�^�_ڃ>Uק��Q��W�g�g��^�v{��=^6p@<Kݬ��&s�:�2��::mww��]�v�+��I'L�b/�tSwPF��̰�o���j�(�L�n�OE�+b�#��Avq��# K٤t>�s�Æ�ǳ_{�1�GЊ��.:9��[(2��:d�II�@��v�L���L��qcG��Џ���:�^S�Z�v݊�i, ؀]��˽'fq����B��r�&�A��b�;-��8-�S�� �p.�P�8��B��A�<l_(�������4���1*,�H�����E�b�F���eE�k��5.}fi%�ޝŦ�N�D���N�oq���xN% ���y�����,�C=)�TB=���=�C��u�����mժU�i�\b��՟�6M�{[63����s���ܓ�t9�9����\q����{��#�����ѣ��ۍ�w|�������9�׿��#�uuY��?�Iw��u3N�iŮv��e�'5=݀`�W�W�wU����<g�����Ֆs����z{bQ9�n#�T�o�hu���v��A��Eb����ٗ�C@@б���m���1Ĭ<媷u��n���b�F0����22�݆�,�Y�uU��պ��!@|���d��g��^~���������F"e�RT����!�ڈS�qe�Ef``D:�Ѧv���6`FF����ܳ~�[2���N�׬����W/8���S���~G�c�X��/�\[[7�\m����X}���g�����S~�Bc�}̽�@^E�D�5oA�؆�S"E�}��G]߬{P�rW>:cP�5�j%�zz����r�sN�q�.��o����="��'K�s ��[䪗'B��C0��-
Id���w��Sm3�U�<obQ�$��bQ�'�KK��~4^���R6���H��i0�D��|\�qq=H;!��=����+--���x � �ٖN�8;m�)6�;v:݌~u�].#+���/t�5�3�	&�5lذ�G���Vv�8�f��f����U�>��� _zF�+,*r�\r�uJ��>å�r�J�q�fS��K�%|�������U��8��yn���Z��d�_X�(FE�Ύnߔ�$s�#S���[�f�O,@gJ���P��6Ľ���&�i�Be�:�g�ǂ��}��P	�qm��x�ƌ�2�2]{�O�]�|���/����Z�7�����w�PB����w���O���'�����&�n��y[��4�J�2& L�E\�n���˶y^��u�����Z����ٹ���0fj�+.`F�r���*�_�JJ�O�2���/��?g�u@g�V�~��j�e�����Y���;<�ݮ��3�C+��������B1U��tY�tΕ������� ]`��[,ʈ����:_��8�/��5U���[�q�8��Y ���8�@U�}8@7c9j,�{��(�h��%?,\o�纬L�A��|�$�L� ��;е���}�r�s�>Q��h\��"`�(+�`��Z��0Æ��'�mx�ر���T�I�j=��q���������Ϟu�Yߛ;w��?g��}�o�Vg�o��'�y����'��r��ܴiӬ�	򨵭�R��/_i{;2��@�o�z���0��uZ1�ҁ�\gW�kjn��Qu!5-�e��F���h�+rj�b���is&�+�^2�gިh�L))�&�f.�~	2�X�i��Vfv�5�6b�ɯ��l]�����������:��j�̨�>m�Y���7Ύœ���(0o�őE&��}=+�����U%�n����G���;]z�?|8@OK�-��F�/��e�A,�oRk]�ǵ6�v�����þ�������k� �֭[?�}��_2Q�L�M����=�x�Y��Z�y���Bp�#��U�@Š9�¡ ]Lw��g���LM[�	��J�����Va��� '�`�g ��,yŢ��C�6E�NgL�3+����r)]��($�-�q�%VF,J
Fx�aXC.u��_�Yԉ .ޔ�4�/�?��x�A�e��(���7�Z�I��6�T�B`7r���6�	p�}�8p��.����ݚ����̙3WO�<����$}�뛁����'?}��/��]�����?�\�ݎ�n���.s�/]����ؠy�Z�����&�ų��N?�t�����]ɀ���jf���Cr����4���a��O��m_�O�Q%_��,g�ۤ$# �!�����Y#�EM��n���}�2����J�X�Y���%�"r���I6�����0����x#|?�#�Y�:'��3��rԳ����L�=i��q\���6x�����ݿ4�"��Wz&�6}����QTXb�t?7�������3�MT��g�z�	'��s����1�������68p P��%:�P�X�hq>6�X,���-�~�C׹��0u �e.K]�cx�Dp����4IY�>$�甒�XC@��
����h� ����m.���Ig!�
���i؃noY��m�<�^�|Ѥ�w��5x��x� ͝�
����.�h0N����.��[�����B�3ּ�㐇�p����cA4�ꮧ��Ι[,==��O}�SHJJ��7ğ�����7��3p�7���>��a��������b.#=�\�칵o�7xM}��ܻ�<{:]s�/	{ʴ���K/���}U��&���=�%η9�����]��)Gd2Z�d�����k�z��"zfz��,ih(%�����
k:]}��|j�/���mذ�Y��t_٭����2�Pp,vda['9�>E��1�����aa�#,�<-Pf�G)>t�ع뗿����`�xg���2���
�=݆#�y�9�����J�\a��7�>���O�t�9�Zt��c�Xҫ�.^][[;��`5o�X).w��{��k�65H�Z�an�����O	c� u��b�q�8����+@��ħ�%�i��=��b�b�����f�$�,Z��� ]�zh��9�OYC揔2��CY"��DEZ��<O���؜�[~�$8��&*a����XzJD�����Qf�^c��N������a���
 y^n.�ZJJJ�w����[RR����U1�w������7��'�x��;8ڟ���=��MM��XJ��[��t+W�v۷�p�wl�]¨VY��a#�w7�p�5-��[����wt����٣ :�4��/>oUܼ��K+�(A��8lͺ��,��"�h*1V,�D��ό���m��wz�QV����cܸqc,?�f3��3��'���;c��"NSr�Ž�р�7�}��JIbn=7��?�{���{�cS#.�{��A�ˌw��������r��.?/w���s�{晳���+� :�Z�f�?TT�MU�::���\��|p/��n��*d��,��$��l.Y_�W��.�@����a��.�>�O,��@ѷ LtŹ�J�c��j�B"P�e*@�?L����/tE'�<!��d����Ƒ�P�zT_b#�$�N1�D=���2O��a�k��o=/]C�Z�|шx&C�`��,��-X�h�l�����'N�x�3��K7C���f��q��?n����g����\�w�u�w�F�j���z���ʽFH[����j��pKW�0x��|w�7���RW�o�+..�~�]�Fp�����-+'=խX�̘�_�r�u�,�=-�
xۺ;�m�s�ou�d�y�}�y�`��9��<�n�Pj���^zɭ]�>��;v���q�����k]X�*\�LD&�6����#8��K�����s�K��S�C��g7e�5�>�����e�4�)�����kO�>��/<o��X{�����W�n݆��f�G� X��=Y»�=�*��d ��p�y�L4�D��,tGy'�{H!p�:�)Rd�j�
�<�<�v����-ND�fjj<��{d~�(�W�/0�����H��}�H�GƋ�k+-�q�����z�I'��1s����@o��%G�����l�A�pӬ} YR��z'bݞ����`�ӦM����|��|��9��Gc#���o�^g���>��?��s�W��1@��/~��
�	�%�u�w��z��^��b���c�.t�edZ�}����X��u�.�,�(MU�N�a���xD�"R���P��*ۅ=_Q�ۼ���
��+�E���X��͞\-c�߸���r�1g�ǽ��5��!�1Bq��]{*��PX�|`NM�H�=>E��Ð�|eP��ȿ���IY����7^������I���l`Tp&�2Pp�z����xS��PaAA�+-+>0z�ȏ_u��8Zk�:|��W��սτu{�M(�n9���Q^��:��;[�Q�S�'-�c(����#!�	��X�zi�,B�SD<)<\^���f9�9�;��.��>d��3����pzx�!��R�s�{��T BY ��=��v�|�	�)Shb����&Y�T�$*A;�C�K���?���h����@��3~�z�z�������S����)'L�ʔ)}�Ǐ��;���<��s'|�k_{}Ϟ=�Y����4X֖���l�7�� ���Kn������w��W��|z��yό���'��Z�q����;��Ns�rl�R�TŤ��Y+Ҩ�& �l��S�.)هT9rU����C9hn� �,��żz�J�/��0yn��,�����8PD�/\��w��b�.�b|*�MN��;z_�\�����L��/����p�lNM�l�^?%%M���P��w�DY���t�Y�v���l�C�?z���<x4�1�-[�L\�n���F�%�	3Wl7L��]�X L %8�̘߱L(���E���փ�gR����O]�d���r_'Z�d
)��y]EB��������'W������d᪅�b�_���9&�Z�~�J��#ҡ>�>�����g	pl{��7�\��y�)����CN�N�bC ��R_������+�E�٘6 1G����1k�y_�2et�M	�w�����b)���]WWW7��I���|��'ԇ�[=hh�RȫV�qo�����XO�۵c�!����kV1}����V��]��þ����.3j
ȡ(�ˁ�'M�����q��jv�T~����MX�F���\B�� W����?3�*ť�&Y3��N<ٍ�y�!{�<�
69/j���Mny��RDi�J7�jJ��&�{J
��*_�zE���g��>�b1��*�a�0���S)�f���22�*&N8���\y����;���`_yeѓ�D�mk���������� i=x3�FR�pw(�[�!&t`v�x�[LwY�r�y�+}6&��9sQ��V���nbL��aH�S�ߕ��fPIJJhy�k����%.e��.nUT��RlZZ�}�޶�(�j�-v*�'et62�B
A)cAÎ��8^��}q߰��ǜ��n    IDAT���L��J(���FW;��қ>��OL�;����-���b��჏�X�� ��s7}ዶ��A�TK ����x)0�a�zWXD�6�s�6W��sC�ug�}��%���Z���Iu�^�8H�B~����g��V���!�=d�0�d�)��6�.Hs��&r/tS�:��800P8ׁ���.t-;�̳\mm�[�l���=_(߬yZ�2&d�p/�(���1oFZ�,ꢆR��\��?4b�b�	Eè�g��Q���g�xyJT���,-)\z�̩�7{�1��s@߶m��U�V�nj��MZ�}���A��c��ܰ�CK !6��� _�K�Y�G��\�e�����4��������#e��#]����`x�9�XF���2a��g�G�T������V�j�k� �L �/##�bG4"�ER��͸�O��'��;=%��f�Ʉ��!#���z��=�z��=QƔ��NKkilj������B���D����7���<��רH���}�]|٥�pKG�)����JsS�Y�;v�Z�����޹ü�4� �8�L׿�āV�����.��j����Q^�����/����{�G#W�D� ʀ�=�\J�j��Fr�ZQ;��O�����7��v��n�i�o\�[�ꢚ\�y

��J'�f���9�_�~6�>�o��8�N�����2c'g�'?���	Y?������8�0�srj���G��0`P�'�8��3N:�U�<��$������~cav�:�Xnf%v{��?<���o&ʻ�S��fgB��@�'�	�墖��x�X�[�VBv���P�`b��u�+���DR���p�P�J�Zb{���X��{9T=T&t���b���s���.(��'ry�>(o�gc����f�!�����q�۾��6�6��MsI��C�4��_G�k�;7+�?�|zL�;f̿��?�k�@���o��g������~���P����ns�9�uvt�Xčٷ�&j?�%��6o��S�݁�z�g�N��r�����'Nq�G���9�Q �i�ӳ�t�p��d��ެ�ڼ'/ r��2��Dmz�۴i��u����&�#�Y�v~B�!��S�N5˚x=�W7X�K�"՚��M�����<;@M�:�mQ-ƣ4dd���Ҍ�3�p!G���ᑰ#���"��@�s.��I��f����sr�+F����pݝ�z��U ���b��UkV���+�^����
IrD��f�s�-ƒ�πD��9~(���)�i��V��q8@7�"��/t����� �O�=#^��TX�P1t��U�T���l����YD
Q����q^�M|1�qo(A��7�a�P�x��C�id�mnvn<�.wcPQ��]࡮G��s��+�I9Ĉ��C6�ќ윻�8��/�����zc���o�f���:����CO��O߬����E}��w��F��Фds�S�έ�w��c)]ٹ�n�>W�{����q-M>����'�8���G�e�h<y��m��iDP���1k��R�4I�.b%%&?�9ⷌ�<c��JZ�'�L^Z���L�v*�!�9V2&;��������L�������=�Z�����������������y΋�W^�sA��������9/� �����!桽�%�.+?���s����>�l��Ə��\����*�΍,_��[�l�YS�O �ni��x\��KdM��K��Sp�Y��9�BO�5�I�˝�����"4��ǅe���(K=�x\��[@�aO�S�?�$�7�$�&��w�����Sd8��w8R��DD%P5�0Ġ1�ޅ�S �=�:1�wД���F,T�|�>�D�~�آ�B� ��I1o�K���>�H�U��qg�o�@��3a}jJx_̏<.ֳ����k_��W��� }�蛁��X�t���k߸��/_�l�҉x��?x@!���.z��k��������a�WV�����l�s�vk�˽�@�k�An��i:�q}��h� ���X�ȀX~6
8������S���\R�{"����g�Q�- ��VH&ó�q_�{�Ve���:�\]}����5�~��B�]�x��h����)xs|)Y�X�[�nw�>���:�T�T��)7�tFH�,���[7�d�a����C�c��O����<��V=n���wWT�k�~]�����CDZ�wQ�3X�,�ij�q�Ԧ4ώ��YK;T_t~�1tY�!�xz��?o��.B���}�g?&��뷴UY�!�]����9����Ʀ�c�t�� �//�w%�����8��E�/�B7{�l#�d�eX̌��3�y���yBsKt��Z���\C�<�w��_�쇮ή?�q���x�Wn=���}3�79�?��{�l�񅍛6�߱}{��Mo��;�7�w��X[b���:�4k�2r����?`�����6m��(�u�f���d@��p�ڑ�|�)�tG[�����벲2\Fv��s@�֡tDD@C��u�D>�>q���t,t�� U:���4%=9b��1lp����[���q�����յ��С�ݤ���|*5�=����}EJ�g�I��Wr#���3ϸ��:�iՌ�4��ק+*��}!/!�b�e�b�ɲ��J��2i���͛�믽��j�΍�رc�M[﫩�$��˗��C�
��7��o�,�U�Ǭ�$��	 �|'$��R�G����{�t�t���Х�X��z�����6�0]���}���b�!�]����^�� ]��a�=���U���E���:h�#R�
�"΃��ݝ�VT�Z�#G�r��k\gw�+,(p�����������_9����~�T��� �w��͹s��,��sϹ��6��f3�4�4���⽗]r�ԩSk�ڛ��z}3�ט�e�6oܸ��;v����=UU��X�UU{��!{���͕�y�Q���ӑ-�p���1���C��eu��n�ڵ��Y��uY��W6p��<t�>b����m-�4+���ͱ��a�M�t�� �:�I,j�
p�d���n���n9���z��e�x/]Ό�V\b�7-F���5��zb1c�|�EG�<u��=��nFW�X�{
�����C�9���֒��YVܧ)'x�Bh�7󔖜�
��s��fd��9|��>�~��X���_���ի�ܱk�c����hT]��[��b��4Y ;w���xZ;�EbZb���b�����&�F�⻤	�C�Ana��@Z���~�)�	S׼�{��Ј�.�;5��x�R����;�����:�E�iXP������<TDt�Ư��!�����W�{�d�
����<�Јq������^~�!�j�JWXPd�d���w^4������?�_�đaC��5W^as�|`5� D
7���c�Gq1�X,�fʴ���\����F�n��X�bàז���m۷_S�w����x�usT�$T���ba~v��]cc��v��_S�ea�o0%��!w^[������UZ(���?a�5o=f�����g�g���c�M��ʴ�S{uUuu�����F��@ 	���0�ˢ��*��������7�:�茊� �"����Ⱦt��}��ںk���y�{*E� ٪~��u�u��sO�s�wy��a��7�d;�^|^9�6��:��]6�;�9����olN�	�r;�� $d���s��A3& 5�����gj`P�H����������Yg�����^7j�q<��CYe�ڻ�S����X<��>��.�{�`g	�Ţ
]�t/�ݪ�R������I3�޻|�����s�n���:�}���o۶��D*i
��Xʦ'_��g��h�r�@�-�)~� %�PVn��� }2�]9q9�;ϝ@]n���:��SZ�T��d@��������n^��u��t-����W.����s�m�����5��#�6���g6r���MD��`Jg���VK�Y���vo��L6��p�����B��l�c61%���P��5c�����<`�B��\U@zҍ)���~�s�n5m��vR�r���ʧ�Z��.X���,����8�f��W�Oݸe�gv��u�,� o4Dg�8:@�8=N�_�4Ia�'�y�9���""�ƻS�^�o��U��v�k*4P~������mS����5}��#�^EL�� ��}��H��μ��_�Z�({j�s"���6s�T6Q���6��l���U4 ����n���Z[����,�����tG�w��G�� �����t��"�y`| J�=i㖭*
3�h6"�̯��)���tT� �S.��zP�f�T�?u�ɳ���/�~4<CG�q�[�l�e���c3z
�]����� u���rC��`��*7��0���סrm�ib\.��d.[�䵵�[���&y�X($�u�]��֡�90��1^,]��>��:�S+��[��������6I[V���M�}9�6FN �p��׫��J��O�TQ�,:��0����PV���P�SS����Im�nȃ�\Gc �У��|�A5:���S���|��ʪ���_��ݣa��ǐ��w:���c�vl���������X1¼�u�֛��C�I1l���*-����S
9�P(��aɝǢqz��B*����P�wlP��$��O�9\��kԴ�'�ٳNV6��AdB�S��H�-pr�rрV�_z��@9��Й��dh��x_�n�ڽ}�tr�(�V�������St����ó_�p��$S�ȸ��w��0 #�r�)YQGF!4����C�V��1Qŋ��T0�z��k��<-h��� !}YRR�l[{�}�_}������0�;b�����踣����cc|�0�:ā�8��I�b�{���풮8�\���Cמ��O���]�\����\��ץ�N�@gx����\@G���k��J��$����ٮ�ݹ =����s����iCg��e��iC��m��X��w��  �I�ۤ
�|�� �]t���6�9g��=�?��B!�C�s9}�4���.��w�{?�}0ۯ]�V՚Ȭu��1A졫�[UVא���#�F �)�~飗_�Ϟ���?��$��4۶m�lں�#ol�������~��mx<�]w:M�]��Gk���f������wC���%[�3���E��]�u �۶��z��GGot�w�!xͭ�S���NWvg:��0�mN׭�@$�_]�Jڝ�E�9{V��͌�Θ�Nc�s�^3�v����_܇�������5sDQg���C�1��8���������w�44��;v�`�{+�� 6��S�V��K �ƺ�ژT��x�0�1uj��o�������:��u�n�����D[B4�b%a--`�����KQq(s�Ӳ���t�р>9���k��7밻>>�D�o�xPu���K����{���Z�Y5<"D8=�ɀ>9���?�	uZ�힣��O>N�[�� cӠ�C:�|Tڐ�=�ܥd�VV�q�B��7�<��s��G��{���������COew���Zv8J���� ��>,F�X��w���(peU��1X�y���;/�����_��x�O���w5�7o�X���O�ۻ����و6�j�P$�gXW{��I�'��O���x7K������/]��U4Bq�u��CA���tسF>�|/��J8ة���JX�L-).SM�S��3p�� �*|":@/F��}�B�wݚ5ܫ�w:P;�b��;���&����Ǐ�3 t�q�ϔ��G���N=E͚5K�'�L��c�����,aZ�����6��,GC: D<���o���,l���$e�Ra�J��oQ�U��.\WS]�ٳ��a�ܹ�]��]}���G�qk[�l���@���~�y �����|a�A� $�n�� zj4k@���sN����k�S{������`�	fxH5ю`9�C��dR�G�C��i�G�k�"%d�c��(������ǯk�ss�޺�ɆΧ�=7
�Ǯ�K2��f�d.2�`��u��6;�_�ǯ(dC�� �}�L���6�ꪫ���XTx�9ތ��H�@f���P?���L)s	Ƭ�t̘1CCc����;����P���x�3�z���W�o���ݻ.m���q0L�D0x�Xp`�,S��g�U9 t�@����/�@}�;�&��G�|�AHED�������bA���k^S��*8��4�34�1�i3f�3�<S�.a���0�.-f�/7�t7���@04�6��N`�8Y�=20(��$�@�� ��@��P����j�)'�C��}�ݧ����P9x���|��>B�؃ ���_��C�G�� �h�"�aRV�����@z=�������ƺ���,Y"�b���Q蘟�۷_�u����!��_��`F��&��ॵ���z����:��jcdhF�oR���<t�:��R3�)�KҨ�ֹ)�CG^W��������ZI���: 	� ��+o��U=�'v���A;�`ІK���Qbf4���ux}"��"B}*ƽ��el΀J�s�I�ie�B����ֹ���[n���5���\y���>�ѱ��1��M0���1c7���W^y�i&�騵����!?��iVm�а~��/�ر��@0\	��@���a �8���JC�l�,-Q:g��X���?`����!:Dh�s�0�z�B�Rj�v�Z�I��Dt��v�51����鳘J�c�`�c\���8r�>a�u���A_t�c/p�HFC_p�����N2� ��4��K�&ϝs*C���a��+*�h8��JX]ba����	���]�v�{�ޏ�X��$W��UJ��
�'*+�W�4���e��~���4G��n�ع��ν������@#�K��C��[��Ń�����aP���: 0��C�q�b�ū,�{���v�C�=t�]���"��t�pi�C�yr]?\Pd�Æ����9'{�����s�r�(ě���@���?� ,�q�;87X�u)Q��o,�K.�0۹H+��CO�U��!�"�������Z���o���	�5�&6C7%�d����1�LP����x�G/�����n��?.?�����ƶ�[6n˖�W�����G�膚pY�IewX��c} ����poHnV%ֱ��2e�I�D2�>�;�5�\�F�d3��:5�vu85�A��ʕ+��МE���"cX�0 x�mSչ��&@�~
*� O�[��1b�i�����.�tPe3�gΜ�����%<��j�PHq�?*�4��: �����ٳ��={��l|e���	"��>s�'��1����,�q� �jw�T���}��r����>���z�y睷��|>�sU�����윶{��Gzz{g��}G"$���z(� h��\���<�`j@פ8]���T���z��ϩ�q:t�P�^��Ҥ8���x��e]Fޟ�JQb/�X{�o��r=h=&��I.��֩��C���� �����5�F�7��*Eb
�ܘ��i������.�H͝;'�Mh�}��С����V�B�����j<�;�\!�&�87 9�"qH&Uyy)S3���&��y�����Շ������ f`���ͫ׬���{/�W�G�,1����PU�U\W���l"��g��g_?�������&X1r���׿��lm9B�Z��zp����.�ݻk'SWC�䱉ו��UP����G-���K��l�˝�4x1��j�+�)oݸ��1��	.\����!�W^�����=�5���H��ɝJ�$��¿y8s�|z��w�����"Hc��#"	�`��c(?!b6:l���Tà�z
�ʜI���Ҏ����O�:�?.\�?����1����e�v�y�Pw��#���� e���J��� ���A��,HT���`rN.���R<����A�=�a��⛛.X�,߲۳JrZO�)2d    IDAT��V-^x8��G2��'?`oE���ssޓ�߹��5|�����9-d��i��0Q���B��P�ق�s�yl
��jM�|�M_|���75�L�r�\�0��=<ux
���~%M��>��;fb1�_�{�c�k�see9�[��/**�x\3���ñ�A����f`͚5�^]�q����/��ԣ�<����`�b_(/�P%%�*4b�
�.}k���o��c�Iȸ����E�=_���u�ɔx%�G�������b��8�.�ۺi#����ZX{���W���b�9�,!�c"��5']�Cڊ*� t��S*�P?zv`����S����O�?ǈ�D(L������}���d$r@Ǿ�}{�9����X���3(o�g_RV��b�W�4d^�
�~� �	�C���v���J�������ϗ^z�\���uT:浿������O]]]7��}*���`!�mV�][��ҬV�Q{��4�a &���N4#��1��w�k(h@ǃ�^����=t�|�l,y�*���.Ӄ��e^�p5c��B�F���s=�\��������.s��l� J$	�x���3�`��4A��D��������.\��3�8�3���-N��_��b���c�E��щ+�dX���!^�9�)(b3B�y``�L*�F�������--Mw�o��??��^��رi��;�o�X��P%@5��2��=xn�kj��6>�gJ |����o"�^� u�7������ƽ�R�O�K��18'Hp�1�A��3���� ��c����7�ۡ4zA��6�g��X��&'r�(7�Ⱦ�\]e5�e�6o&	�g0, ������y��<��ȶ�%2i�[��I!�  �keM��9`�?�����-��0Ƚ�}O���	O�/�k�UP�;��VW[�pKˬ��,9�䢏Z@���c�;;;����w�K�F�x�������%��: =K21�st��OR�m��b���9f���f �̥=���z� ����u���6@V��L�����o�k�Y{��r�����5��\����gث��O�)�� ��Nw0!���f��:��9�2gΜ�fΜ);P�+��؇��or:]_	�B-h��V4�)�^���t�%�n�"EHN�^Ū	�7{�L��``##��S����k�d�?����f`͚�֯�;w�o`���L,N�mL NEE#o�`὞�j�c/�{�#Ԯ+^���E�X���5u�eU���YQ B� d�<��`�ݎ�Hip�t�	X�(S���~�P��8��Ş7�Z��L5M�P@�8/�g��@@G�l�֭��L��M,k�����^��
��a��\���0����-R���p��V��:�ܥ,{����'r��;���x��?Rw��d�K�f��������[Z����q�t,����;�7�u�֏�ڵ�'�㑆�o����F��"�o�9 XBPϪ���\L.�kp���uNf��[W�������%�q۬���*�h���1:O��a�#��
���֥�d�}�/�팓���8��D.�Jˬ"���g����f:(aA����鱳�^��˖�3�U��ߐΘ~�F�����aq�����á����Bhn�����=�ݳ�eoؼ�-[�|ii�555יL&	��_�x�g`uGG�Ƶ��ر�����]x�X� jD]��U�<���-�*�=XjM���P�2����!��k�JJ���u����ĸ
�'���x�݉	�	�i �ڥ%�<wW����l��H	鸵����ݻx<�7�?�Yj޼�*���(C�联�£ր�j�]۶�QnHĢU/��۲v��,����n���G:#�I7���>��-��7��zG���;�S����+/-��|[�KK�z��_.�7��}~������ۿ���{��`W��x �B��W9mA�ߥ|M���{ՌO ���Q�1������u}N>@Q�p����s:��c�hA\�R�l�#!�`� g@���o��52�
�1�\�_{��{o��ى\�ɀ�=t-���Pv��u7���l�mS^��G�͛���������߂���!c	����.��H����hi���c���H��T�����mmm_1�L���Q���:Fg`�֭��n�u�[ol�����r.�R#w�網��@����8�i��,�� �._V˛�d\�ٰn�?���;��.��nR��U V��1�JF�$�\�T�`�y��ھM:�eRg���}�ڵk'ذ�������FÁ��IIY�v� �a��O|ώ��"7O��f��-*� ��mo�S7�Ҝ'��@��RR���c�^		������N�=���}���NH5�x�sN9��C۽���S[�����K_?F��<�c�q�;w�,�����7~v|<J� ����;�K6�&]�xLڲ"��2+�\�ԡ0��p<Xx�q1�[ :��u�Wz��o8/<�(U�k8���x?��q�������s��71e�9�|�Ѯ��DhȨ��p�W�2{����z������|��o�[��K�d� s��+�(��a��/�Q�b����q�a�p8�/Oij����b��1��9�3�;7v�ֿ�ʭ7o�ˑa+@�������8�������� 84<ȵ=���g��h�%��S�ZN;%��e͹ɬ�����3���aF�F�ա��{p`�@��E��n�6qq����E�ͤ�ْ���fU[]�֯_G���U�D@_t�5s�,5�F �n�Rn�V��n--�zݷk�R��ø
�΂�J��PII�����$�`����`�����h��W ��o����v���S��N����kn�?�<�D}z�)@�_�+��rņ?��b��s�uѧW@k\{���>��F%����'{�B.�k�|�'��5�GK��}� X�\��".ZJ�C��������A��PE���P�AJ�&�rs����	5�����������&�
��2�
.z� 
�T�x�����ŋ��׋/�x���`��C�d2��і6P?��<��4��)t�s���J�8eʔo����|�ǔ?_~v��Q�چ�^߰�־����Ƃj,P�h�%Y�2=�W�U�u�\�X���Q�g��A�yR�-VJ��L����x"��1�J'	�� ��Ca�O}��R��X�F�j1������!�\���u�+.bXzxp�e��q񜓉U�`Ɵ�GԮ�;Ծ}{��ȡ{�>u�%�����jhx��s�h�u被a�> ����V :��Yy�<�c-��ױa=y8V��4�R�G�����f���t[�u��?�И
��'���3��pho����o�ԧN�'��t|Y�7o��z��G��Ҫ����^"����I*!Y��ix�Q��>EE.�\�;Hs��\�9[,�D\�r�΍�$�r"7��t��h�@�{!wX���Z���d��N������:������d '��"MR`�P��j�}��W��h���1c�.<��Fs||�6~����/FGG�����8M�j�y<��>��>��)��7z�.��}p3�m�6���;�ݸq�]=�}��PC��u�g�$\�+)V>o�S 0��7[�C[��B�u9�g	����"��9~V�A2�Z�����ޣZ[��ట���ݫ�Y�' ?�5��oN��"�
)������i�$��PSgL%)ar]"�H��N�������;�χ���J!�Ŭ�ҰD�Vש��Z�e�j�3O�>ᘸ\NUW_�����AG�_�5�骪
)IMHc.��sf���_����Ë�=�Rɤ���(�M�dQ��
���濹��;���������,�cZ���׶r���l�i�棭T�Õh	�Y�f�O�ǣYb �,yе��C^P#?�v�.P"R��M�E+�p\��fv�3�X������E�t��!<��r��g � ]�g��o�L��^,O1�}9o�Ii�#$����<w�����k���a�hV�B��2�����������x�{<�.�k�d2���G��Ϗ���G��E:��ߞޞ�#~��k�\�,�#����+o��%! �C����>�Ak�(��XV����]�*>��5��,$r
����3�!��,\���󪶶^��62<F���@��b��Y�dbq��^�U���h�`HBډ�\�0� f:�xf��`�����W~���9��bqQڔ����,sjll��gǦ�j�˫�(�(��RR�U�;6����PQ�s�R�ƭ�*˄e
)��!w��B�u����_W����ط����q��p�:묳��ϻ��k�y�D}i@Ǘ�aÆ�C�=2�����CP����|#.�)�K�_6X�X8��iK�>�[�F����FnY�=>�k�����(X�X�8^����&�!�%�w�r�:lY����1iŦ��Eй9���霸�_\mY��pl�������g�zٲe'�����9O�\9�+k���ۿlx�o�,e�X/X��X�b�c�`?�"�~����t~[x,��4H�0̱>�I�5k-rz�6����ج~Ww7[û���Wj���~���T��J��1��m�d����6<��n	��H�J��V+��>r�F�!D@���C�})��N;�Q�آ��EjӦ-�?���ae��ϓQ�슧����s���yQ��?�l�� t�o�K�/�
x�8$_�0��o۲U���(�IFJN=����.���%K��k������/���ӷo����n�NĭT�V;�4�3䎞�hz`�^Gh^�;=`еg<�C�-_#Ъ7���x���Z���
p�c�#珅��&�3��DN.'�]��5���Z*$=~F�={=^}��s�Mfu8�O��~ߒE�6ͭ��E����k�x��^[��ˇ�{.�=0��'9�j'�b��+����Ǌc � Bԓ�6��3 ��&\�ʱ�t�G���xSq�.,T�p�&�\�3���^) x��.澑7G��v�� ������ JƹD� �0 P�.i�$�ǘ0V�������k�R���@�e���A��y�p?õq��(��0XRɘ�(+U�m�T��D��Ժ�8_m�|�YW��E�_�5�& �t;%r�JJ*�(��c�6m%_ۧ��O<�ƍ���;vJj��q _x�E���_��5G����� t=e۶m�����``��(�b�2�@�lt2%C�n��tQkZ{ʹ��ba�|�����c��E.)�Hq�{r�1ԲH>���gIn<��8���x���k�������v��K�K�p�I��ԧn��p����3p�g`�ʗf��i�Wt����ǋ�4�Hx��*���cF�*����Mޘ�NIu81xi O ���p���C2&퀱O�3a�/���Q��g>�jjꘇ���W���,7C�9C�Q)5C.?\���Eʼ�$`��J�9��1�9	�85�K/Z���z���ķYѐ%��5"
.�W]{�m�4~�81�x����I)�)���Teu������ǟP=�}[uM�jijT��^�:��r4�V�р9���e���1�Q���I3fR8���\=���L�b>��ڭF�F��n!����-u��eK>w��V�'�ȍ�t�[�l��p軁��T ���a�ᑑ���4i�Vz���z������sY�C�Xd�H��`a�$]��f.8Ub1Z�X�"�(�8�	�1�u$7>�u8�.�����N^�b2�66�=4o���.��¡#��寜��#3+^xe��뾴�����GJJ�v�	!��|%��P��#B�RO�O��Ւ'�� ��8#��}���&�=����ᓟ��������vq/��`���P�=L	�$:rs���V�%��8�y���9��F@��|�g0�����Uow���&�5��f�?�����W%%e��?��(Ź�XW�]UU����U�t��^Z��La߃<+��=����<v5�)���� �.�B��Y�c6��7s����� �Y�"�s�vjV��k�[���������#�D=W=� ]O���/ھs���F�
�܁�ԍ�a�RS��E�OH��W��O��yt�O�b�o�'�FpF�V2�s��ᢂu<
r�`����f�����o*[����ʽ���E�M�[�b�q!�{c��33fL��/~��K�����G���w6+^|�i�������v��L�dZ���J$	4�; ��G+�І���ÿ�g kǣ���)��� Z8��&�2Rf4u���pH�O�������c��J�� {���9vLK�e��J�=�R%�p8��\wl����Z�x����h�0����d��(@e���`��}���#�/g��|�h����ˤ�8m���R57�QO~���y���"4�g�Z�a�JƢ�q�~i��,��ө-�!x휠gǴ��3<r�>߹o���:�\��O��3����ͷ�p���ӝ���S�?u���m�c�߹��=��g���a�R�5�`OaM�c����N]n�=�oe"�E�_{�(���3Y��$�`21�0����G tX���uUm����������9���g�(-*���g/��MW]��~<0�s�g�X� ��u�����jhd��t(a:d,�x��_��H;N�3���������~2�u�\�k&�-�p���
 ����&�P�ļ�wuU����+ե�_���A������9w�{����F�oGJ ^�n���E�@�Q�C�d�x���{p,��'"!��a��D�4`qi�*p����^GA�@0dHʊ�U��a3ʨҪ�ԧjj�TCC��?����F����|�Y��sH%IVH���յ�C�,o	ct{��A���̧Nkc3.�ɏ���>��C���t�Oo�7���E���W��:��{o&�1����PW׷��@,X�:J��!C�Aw�`��Rt����s����E�gny��$yv	/��8�7 셅�o����[kS�FFZ{{zo���ySgg���Z��E)]�?��#�c9N��c])�q���?9���,[�l��Y�3�8�g�厎�V�x{Ww�M�p��`������P�<I{� r��%E�K?	QRi��.^'�p>�\ue�b�Kþ�iɩ�􅵏s�t�I��nS�ͭ,G;x�� �(�ب �����#��!@.��G�lRd{k�8x��+�>��uR�#� t�ـd�h`<:�27��"��[�N;�tu�e�S� ����N=�\_�	��P˖�UUu��__���/[�����?���ڶ}kv�$�����/��5��a�����b��+qUUU��7�;x�`��`�D<��ok���������R�<֟u=���������ع��=ݟ��Ce)@��ՠ�41�K��RIdw -	�sXg�vfCJEt����҆Z\"KI�6��h�o��Y�f�����M�CV<�܂կ���ݻw��E�#�a����b���'�;*�L'���f�:�{K,X�g�/K4�v6n��{���o������LagK4��l�����]� �0�Y���G�Z�X��IIi$2��'x�Ñ=������Y� ��v��v �!W�y�>��`��x�40G� `��v�$�����K?uDqo���sh' {�� Rx�Y�x*���_EU5��ŋ��s�,ejr,4���W�u�; g���B��4���
����B�W��z�e��u��t���1�~���F�q�3��aap��E������0<wΜ���w��a�%aM���Νx��ŉp�	��ݵk�ɛ7o�����s��2�`���l�o�tEb�Lx��Aư���/]7a�o<��L��h��������kjj^����\���l���Hx�F��ai�!׹u�T7z�8���]w�_��OO�U��Ƿ����N�y��ޜ�N    IDATޞ;Siu:RX����8�"��1�7�<\����=�(z�跍���\��6ڈ
G�,[3�7 -e��</����+����ݍR�����а
���i�
o®(���E�	ֿtT���!���ҩX��q � �!��1C�@-ײ(���1�Ta�WM�q����+��Уzz�X.'Q����ŢF��M�����V�7֩�G=���ʔ6�.��_|A��v���{,��O� W ez�dL&#Z\Tȿ777��O>Y�:��.?�����w6'$�cj���߱c׽c� �&a!�>�xxu^=7̭�U��9�vCz��E���Bʾ�>:gΜ�>}��w�u�Q�<��ikּ��=���Z�V���a��\II�ֲ���-[���s�=��9���o3�����6m�t{*�Z �����p �rW l�5t����q���? M�*/)e������:Į��a�GCƤb	!y�<�N��n��FzȨ[?p�K�ر����x"�H �����������|BŢǾ��#g��H�h�rX{��1f����ziP`��Ϡ�m���h$ېzX�e�9sOˆڇ�F��X��$b�G�=,�mh�Wť%h�Ʋ�D4��~ׁN�v��nA'�q���-���1@�{ƈW�CT-O>y�3q���?m֖��y����t=�h��w��;:;;o����x�u�IK�X�pן�"�av(%A�$�������_����2e�����=��cS6l�xa(<+�zLs����ZCk�S�����$�s/���g�����~�����o��@��X� s��07^`[#�\9n�k0ʑ#GK�hL�;�H�6 ���W�4��p��lD����q�CEƥ�2���I3g�˯�B�r�:
 ���ܯ����!~6B8�㪪�ar�:*�k�C�0L��[�#l4і�d�DV�0xa<EE�����>՜!��m�'�댅�E]��4}�u��cO��p�1��|\U�����V��ܤNu`�Ar ��A}{g�>e6r��t����T���$3�b@$��}�(�?��ST]]��O}��y��w�rNx@�S�g�oWW�����vhh�D"��{��ߚ�~8�n�Ǌ��:KKK_�������ٔ�_��0d~��<�����=��=����SUoUwc�#�Q�Б���[<e���%ϭH����Q0c3��Ji�58�w���X�QO���_��-X�����ܵ�yy]N��]�HJ������MB�pݗB_7�2��J��5A��w4UaM�ۓ%�H=�t�������ڦ>��+UYy����eɜ��ƹ�1�!�tQk��SmӦ����H]�j���{�xϯ�k<Je7�2Mi�+*����j:������o�������⒇���q�~&�o��oڴ���wx�����t:}r4�H$�0��f˄�fu�
��\k��Z_u�\�3gΔ$V�����|`3�aÆ�G}�{�����2W�&bj,��)¾��o�g ����QK/URj	vC����V���Fkc��f--��$��KK��ї/�@9�j���PW�ڳo/	p,+"��0�q��K��!d� ��3rx� ����jg:�"՚P��������qm��bwp��b�
v��#ea�g k:�`d��/VS�N�"\(�v<dX#�t��CB6�TE�B��֪Z�4���5��m[�ӳN'�l�r�s?�I���x�`�LJ� ���nS6���E�ڧ���?��Y��Η���Ք�w8Yȹ˺6�Fl�����|h3�v�|��v���"�ȩ �����R*�Ȓϐ3F��fx� ;��@o���G	�"��PN��s=Ɇ�u�:�D�p�p������T˗/���k���Y6a�q���*F��c� Tx��]��,<a�2pFBBD��J�"�Y`W��@�R9�9Ș�g�9�!�*V<C��qL�"GҜJQc^H�V�`��j�G��]݇�]<k��D�%r�`GK�ӧ���F�+/U^ߨz��iD��/�2�|̝�l~�	��a�(v�COv��p�Qimnd�zue�o��k?��8�PЏ�/2�8^gࡇ~���կ�;11�����c♂�`-++������Tc�Y���� $h��+*a)�%e�P�i���h9g�S��J)�h�iemm5�㋗,UG��;w�&s�<�Wx��j�� hžR��dUja3�H�%��D���0���[������Zh΂��+Z����1�U���7" ��{���,p�m��|�*���Ą�>�u�G.�!T��D�/��x��HXJsM�UϞ5��X�lS�䊧Tq�������%�%���x�N����:� 0w�����'�e�JMk�Bm����K.�t���3�A�W�?��͟7?���f�x���g��N4��4O:ᑎ��JE��Png���^�mi����sd<D0� Hv{��g����\t�f�CA^�.0C�Ye�����C���C$�����g�P<� ,�*�y��q���#*	2����U��a��9 ��w�OX�Z�mXS���$�����a4 |?<=� �%k�(���#"P��ˮR%eU��E����lK�i��ᅾ�0J���Vש��U�v�R7oRՕU�x����A�!�DB��h�!�7�B�ۣ
�E��,��@?y�UZ��w����<��?�T�g=|���~�~q�a�g�x��իWW��cO|mph�
��^�<1�" 4� @8�ZI)C�� �69f�����m69>��- \�RN��D^���=��1��#?��9<���HP�%���Ҵx� ~��n��������N�x*�(����56:�h"�z�t򞴠�v��[�x��Q�t0�� ����K������t2��Uss�Zr�y���U��Q�H{`��z d���E/��8H|hiZYQ���Z��U�7X�+W>�cc���Y9`4c�`�#�ێ)��P��V0=@�zZ�Z՜ٳTqq�n�������y_y@� g7���g��@oo����[�����v�}@l4�>�F/�)� N /�(���HzK�$��tf�_o��4e2�[��IQ1@�k fP,�G�7��1�Շ�~�����8=��ȑ#7��n <�� J& 4��$c*	�@@z����: �PT����k�'D\�Q������2�+*�q�q�-�����{D��
�S_�!�9��)�oX��׹���G�V����F"�Q�E566���OimV[�تvlߥ*k�վ�{�֭[USc=� ����Ţ�T��0j�U��t ��[d������Qӧ�g�ڛϹ���O�6��x�L:0��u����@~޷��o~��+���X,:�� h �ւ@����
8�{e�v<ʰ������QS܆�2�D/Z�wiat��rʚ����A`;����0p�`8L%I�#-V���xɨ��::r�1�
�ц`@�f�aܟ�[��8	mF����i���aw����e
��@w۶mj�����f;X%���-�1ƥK�R#�1CãbLR�f佡�ik-���y�$���.+|�e��Jf���V�T3fL#�wtt�E/u�&(�����ܽ�2v�ܘ̪��\�67m��#KNokk��o�	t�<��@_v�V�3p���K/����������6��� !l ֞"r� �Ҋr
@�S�zz��?�VxÔj�x(`��| 4��P�D��J���𫪩�w��u�ǆ�����1v%�z�`��=b` `�t���W�Re��Ġ)?���!�2��(�`݀u���È �#'��b��gL�I�A�*��L��F3��ޞ�\lqq�&ыA��Yg���4���]j,(Z�Z!�eԺ�J��;�}mu%�o�@l��5�WS㾩�)�v�Z�60>���.���R��veF3(�M(��N��ӧ~��k������+�����M�Ǚ���l��n�ؼ�%���#�#j4(^"�E0��;#w[['�^x_wK	=���s�7�}ޭ�k�׬�� ,�.�P�`�F����Y��s�� O�` �:Px+-+W%�))�I��@�E�I�z�1��?�B�0T&�Xp�/ΟL����*2c]}��UY�;���TLv�΍�<�Ҳ�l���Y-Zt��X�hp�܈4,C�S�QK��G��j0Z�|�k;S]!p޼yC;w�,G�@����"���U�����"J n��k���{ss��ENY4wn���{\�y@���X~�3��f�w�{|�3+�y0�H/7��=*��0��A�n�қ�^/j�<�FIފ���-s6_�G��p�n��ÿ"�"-Nu2 ��iG،c@X]�jD!2~�<��ںz
��\�.i�%��1):�ln���`��E 袍���2U׿���I1to��Ir�PZ��n`���P��\ 8FF{UU���-$��(��Ϙ�@������d�݂U����
�U���: �R �0,�x�����z}}�Z0��h0`Z�v-��9� �{|��YQB0T@�K�c���hii��O��O���*�)F��Ӑ����g�Ø�5k�<���/w�?���U�m�g]" 4j� ����E8^��n7;�0��skyS�'����&@\k��x ��$ '�F75KV%�l��!�����ut�?�9�Kǣ�@׬yx�8^���T��S �ilhRu�����?$��CO$b�W\D/�zwO�H�67�(�۫zz���?��#`��s\ lPF�H�C7J�{���K��2��Z{��k����k�F�Mm���^?w�֭> 7��jsd[HC���e��D!�*�@Y`�����/\�𤏜sΞ�Y<^��������W~��������g�]q��n�_�.Tc#~*��G*<!��� �� up�O�Y������ �x�/]��`�-A�d��,x��p:F�Y���4�:>.!z��+�&���H�z�|��:���x�!Iav]�FVzT�fZY�P�s�xa� }�լƍ�m�����JJ��aE>1����g �ˁR���[RZL/!{����S�����$��
�	�0Xp>���=y���n8���C�������z�������jY�h�Y4̚������u=}}S��z]�,|�2۬�kD4���y]1񘲚Ӫ��\�4�>z�m���Q���C��1������cc����/�A__�����vl�hɉ���1�O�Z�h���*����ޜ�n*  ��- �uX]{��6w�[ZZr:����Zt�b&% ��������/>� ��B�ZK��Ct�5~H�2|N�@�Fwu�G��ᓳ�F�� ?�%y��Q�$�����m0� w{�<�����,W���̷㚃��d���������8yM����"R��� ���2=����f9{v�z��7�t�-7\��o��w7��?�����ez����
#�B0�(��ysN�8�E�.U[S��^�x�ҥ�^?6��w�y@?z�����3pL����oX��@yy�i (��$�  ]���'��s�T��� 	��� �㥕��i�" ��u{��lΉ�iO���%�N�@Y�T�JJ�0.�S�p/�'cA(�o���ka�G�24ir�@��z������GM]-�V8vF��߻w�:���s�����[h�k?rѳf��� �ȣ��C���N ���~���X�cn��o��Ĝ���h�h`\�x~����̅K�to޼�}�ͷ�:2������>W ��l6)�C� �F�B�3�bͨ��b��X��;?��K���(|Џ�/"?��/3��}O����B�������V� ��D\j�#���XMʬ2�+�VY��N\җ�RTTL Ecx����@�=��V�qj�;t�J�tm7eL���;��0пukU��"mI�6������M������F<  P ��)4@7^�D��X���ԤZ[����)�C<U���W۶na�4 !<rvTSj�cN1W�B��M�9��GΜ��PQ�Ϥ9q��9�R��S7>�w�����P;�R��V7�����s����̑\��k��q��oa�ieL���!��i\閴�چ� ���P�奱3�;����o>^��#yy@?����v~����o]���x
OG�5OeC��H�PYJ�Q�V��IJz�k1��.��$�С�aCY�ts�O�3�P����D�%*yL��4� =�����9ޓ�Ɣ� 2�M��5@j�V��/j�t���񪆆F��Ԣ*�����tT��;w����	Mi��8���{D"���ԩ���;K�B�E.�=4B!�����v̭�����X��n�a��38��g~h�_�����O�|�&���>�{���tڋ9� _nu0�my\�mj�Q�M �ڣ�.C��i��y�Ǐ�ep�n'�Gl������3{��q<����޹sק��j��K�艁l6�axz��T@�Ue�� <��݅�������g��d����qZ`�(<U#,�$�d�=rĸ�n 3�j����U�O9��>@�t|Js�#�9rmD��ܒ�mo��<��E���]56����R�t�T�Uw�!�ʻ�'���.p)���*D�ܤ*��~�GE"jhd��w�G�����b�_XC7�c 5�@��
�.z���4��{�?��s��/�����|��r媆{��W��D�������T2���0��v �I�9�nO��BUWW3�x���h�����������8�g`�ڵ�+V<�Hx����&�H��u r�ײ,��RO*`)<6�³ 9��O��Y�	� ��WP)�h� ��N$Q�F�;�\�q6C���yk!��4y��3r�37Q�M�^�(9vݍ͊��N�ux�`�#* =��`{��.�a�1gh` �bo�Ҧ
�Ū��<��m߾]u8�9��`>�/�OD�E��4�nQn��Q�U���l�������y������q���=�5
�+����6� ~���� ��P��S�|��w���z:.��/~�}��OL�b������(�˭J�JYnW\Z�,&��GB����,&���O�ҭ7_��1� ����Q�e䇒��cmV����=���V��jd e ʪ � %�K��lyl�讕I�	N�%���Q`DS��u� �W*Ʌ%D, �Q�Y9l�,����� ���-)�!^�C�Z���!@� xz�FnB*0�����N�pP�����י�EŐH���a%��p  ye�1��28x�l��ݣ��ߧX҅�y
 �"�3����U����1�ntc!5��{��:��u�]葰�Jq���q.��4;�S�u�����Z�xt�r�UUU���oB?�w�}�'���?���������+�P�����J��?�0��QT2�T��P���l��ʏ.hnn������2y@_�1���X3��dlϿ��[�n�+e�XZ��2F�/���	i����6:��фJ'�<�
 �{�m@�v�L��	�����>���Zh�` :kV�`%�4�����л�8�	{=��ڋ�z�c�M� ��J�ػ�%����c�h�� ����:2�H�Gos:h�h�x�-C( kw8U�Р��<�zz�U��tF9��P�(�	3lq>0@.�r��%��j��[�o8����kY�x<�<nHؖ� ������!u��Ae�;���ӷ|l�̙a��O�Ţ�����Jg�6�"���Ԫ܅E���AU��*����ub4%��ȰJ���nU���B�9�������'O�U���m�?�9�_!?�����W�ٻ�?v�ۻ,�ʨچ�Æ��futx��H�;A�5�nn�K9�NUV��&"܂�e�OM��IP��*�ze�Y[��Y��K@��8�Q
��ˑ��з��C�^�0�EPE��k�+pڦ    IDAT]��P�3[�w��3f�ei	e�I(ܔTY��Q 6���mR��L0E@���R��)�B	ڌ:�u����E.�f�{ AMԺ��;..�����Gh�j�qn��*��̫��k���8�FJA�*-)f�r�0`xa< ��OLl����z�\C[��'_���׾�X2���y�A ��\�UUS��r��t��F6�
��H8��jTue�o���]�W��(��<�%_D~�8f`pp�m������)oQ�J��C��y׍7R����hnbV��bi�RY�
�^5�Hr��^�.A��5�:i�CDP XNG�,�񰊄��)� l�zz�Rw}��s�?趦��1���Yo����o��c�oj^��;@1�е�\q-t!����L �=�7�b�h��z�������趆륓ҏ  �ox٨��`��5~�(+���ʊ*��Q����u���BLC�H���*����:H��Վ��n�t^���/Y���m�����~����z2�-6��UYQ�ꛚUYy���>���N�J���Ŭʋ�{/:�ܳ�ϟ?p,<����~�}c���g�� ��`W��`�`/�=��6���}��!�y��ڽ{�bh}�<vCY��������dZ@�ñde�SX�`��V� O�7���`@F!�#?�+�����7͞&���gx�8�C�X֪o ��DX:��D$פ�`(�i#�W"JkTc+*���_O_/��0�P�l��OY��@�����F�8�L��y1��J�/_%��˹B����=�TZB��c|��|�L{@I����za,�.���n�����ɺ�����c���C1V�P��jaos���j�ŊgaB�"BD� ���*e�$Ԭ��>���~�=���e�~�������?~��h�ώ����p��2���e�F �o����tdh��5�ϊ�n�]9�^e�;DZO<r8�d�9��
J�D�$8�V���Nde_�'���H��'�MHq,C3�pD�����lF��Kt��ȡ�s:�@g: �0$�	�\�\�;��C�� ,���(��|\�"}�ǣF׍E��1��=.M�|����^$U���y�V����&.`��q~��/-��V���@B�CC�A�c�ܹ�}�Kw�D?5���ُ���K��qw2-��O<� 鮺���w��AD{V�(���S�+�ʲRUYQ��W�tg�\��?��3L��<�矉��g���M��|{���_G��x` v�(_��:04H�ſQF �:��-�#���e_Y�**����qF��tR<_ݵl`������AC����n��Pפ7�e�r3���s������.^�h�Y¨ �RB2)�ԏg[���KT֤kZ��o��C͒kGV=�7ntC���o���P@H�mWCh�*0�lRf�԰�|O��\�Ѥ@�Re�<�{�;�Z�ByE)� etkFU__}��3���o�s�	�Y�Rw�������?�Ng�a��B��-�T�e���}�*���
���Ѫx0T���^�k��W^�x�ܹ���Ö?�=�@�����?���c:��������k��{	�ᰄ�Y��HPb%�NP�<cx� r �Q�S�C@���Ч�n����+O'3*
]wH��2jl4 �Q��)2�ɀ5�x�&�͙��f��*�2   ��޺��e�I� �^�#g(YY�^�>z���O'��c�,F��D�/�� A��c~t��`�H(H�R���$;n��M��Ek`�1��і��2�u�4�	�#�D���t&v�v(O�t�õHT�H~C%� 3f�x�꿸��˗/���{�w���7��e2�jE�tp '� hnmS��4Dp�l�2A��#�ح������K/Z�ĉ�b��]����}���8&f`�֭Wo���k(�mڴŐ
�r�D*��k:���,�M�q���S�yUqQ	�u�`U�20 R�m#��%�D|�&<F�mA�
��( j�q�u�}6܍���������`�� �$���*O� GM�#�+V%E^^2��`��DF�_��%��6��t��f6� ���\����u4C����P�׍%�� e6J��{/�(�ọ��%��y�pO8(����=��h�z� �{�s�f���Zw M@�������+.ށ�>��?N����uE:�ib�?)���HfDμ��Q�Dn�0��1ԹG9��̚�Y'����}�����~�2����~~>�X�~�#�w����͛���[��eh����^� r���BlC�W���]2omVK�"�K��<�3��v")En&@���n���e���5>���I
kϑ��I�Y�q. ڀ"<�I	]h������oZ9N�����o�k���$�[��ъ�m���$	�èi�Pm�l4J��B*%o`���0�D�D�!�p,��'"FT"ͺr��{�u s���E���k�.�y:�����~����|s��������?�̦�4�� �L�WT���@�9	���M�06�g��������䲹s�"��}�3��x������>O?��������ݾ}'A ��Na���2ja .�{�� ��������k@�ˍ-���J�:�qiԂ�6�f��a2���N-6{<aL @I��I~��W�+TS3Z���)�=*�gK��B�z��U08F��V#�������ؐ�q����^�w�1 �9x�&&$��\9C�vԔKU@��^�q����PMotTw��lY�6x�Y��C@oh����O�E���T��ꫯ��}߾�8�?�Ïg���Oy�}�8?����v�4�eJ+��U<&�	xP�KĕŔQ>/t�+v���,Y2��X_����~�|S�q�g���c�?���� ������W0�Y'�P{<%;J��'N&T�x��o��YJ3 #TYD����4r���4˨#G=��ۤ�	A�j�<��x h�<X֒���#@�������;�ˆ��CYB�����k�@~��c�$A/�~����Q�����R�`{Tz�:�ow�++��{�&5d�#�`D/��� ���+"�3T���X���;�CI�rTttt�'il�ҥ��ˏ~�c�᾿y`��?�G�Tj
���P�ޤ��U���jUs���qo0��u�AA�v4�1+r$*��g�?�]~��#�؞����	���o:?�|�^�쮡��v�]G�B|bK�xb�F�S���PW*n�AE�<� X����gq��M��ʤ�"�b9�n�<%W�E3�A�Ӥ7��Ή3$ox�҆UYB\K3-@�e��k/�� ��zm��^�&;�� �Ei�X��}�-)t�3B�ӆ	 ��v�}����Վy�:��g� h��KEQ�W΁����hO HCc<�;63r�RG�s�
�B �cN�~4���1zԡpd�ܹ�~������կ�7�W��ϧ-VK�n0C�Z#EPYS��Z��Gٜh�G�ب?[o�9򸤑̼9s>��O���w���|?f ���,�ϑ���xּ���������7��� t226�BA��c�Ē&����a�jI(
|����JǴ���5�k2�.)��A�C�.���G
�@�.#���SFW1\F��X�c�kh$�Ⳑ����1��>\��9v��)�k0On1K�?����G��}g	x�ȍ֮���I�F<da+�\9rӺ�a�low#d�2i�	�ء��(B�0>a�|���D��l6�O�9�������0������y��Gm6����c�0X0��WU�֨��֮C{r�Z�/�C<N����Pn��}�]���q�$��[��Q�������cv��q�ol�96qx��F�"y
O�d=pl���m6�b�9�a94���	.�� T�1�͹�^��Df�
� ܍�;j��疦iO�%J���t�t�u !B� �a�4"7 F
# 6{V��� �` :�]��iv<<d
�$�F	�kB��Fu���]HF>��Z��l���	�}�R���h ^�٤���4 <K�`p�{f}9�	/�g:�I����������v�_޽��'�n�����H�"���}]����S��5�MOPD�](P)���īR��媥��߿|�]��L&Q�ɿ>����:����g�؛���^׶�_���;U�n�) xP:�ŌP7ۆf�c�e}#�E]���R��F#�\��R4M.�� z��	��O�
��Ab@�3��G��_SW�I�P��ٹO���)�ê�Vh�����c�CF䁯4��i����EX���(ۋǒd�Owp;,c�A����\��!x�o�Q�.|xԸ�vS�5��A�{cx�^��%E>:������9�'��a\��݇�p$mni}๧g	ٕ�������z����b^��ͪ��>UR^���Zx��-m8�qI'������7/**T�uO\�|�U."���g ����/���co���{ڶm��k``�:˔�QvQC�]����oIvH���d�1�E٨'�g��fL�Jf��6�i#/� @R5�" \ R���;�����Q�1Q���E�u���T�s4.�g����	���U&z���y�YU%�J�$˒�8��'G�'�1q�@0�z5	�8@?��f-�z	���4d�,��L�q���[�\R�U��u�����ٷ~Wbb��}תUUw��s�s����O�"�2�ސ�ݪ�L=�[\DF���5��x�����I�y�����զ�2�����5Z����R
��(�c���U|��:U��+���''�~<A� K ��ɓ�)O�t�[��k�������߿����-�w�ر_�{=������x�բk���Mm^�į�G��d�9H�Q3ŕ�	�&���7=��[oy�޽{�o���=#VBԙ(g�cǎ]q�ر������:s�JԿ����0K��w9�y��<^FÃ�����F���\P����@����)a �m۶�C��8u�|��&-�� =֥ٟ=8��4r���r 4q�YM��2�B��_��7��8����^��:Q�s@�؈{jd	���σ�)��ξz)��\rh��4���[��S�\O	,�\��ih��y�:��p��\�K�W�������Ýwޙ��O��_...��j�"� (�{�����q32���̑����Y�J-P@c�R6�r�ƒ���l�|��^��sgu�ſ/J��"}�"�G�H�R����������R1OT��b�>�m[I�c���:Q�-6I��K��6!5��%@D���Om>A�&�=;7M-9��p-�F����In@r�u�����>嶭O��\�Uݕ�H�W"�qm��Υ`aA����ͪV��JD>:ǁ��y������j���Ճ��vۄ��3�4������Q���@kS\'�.�j�D���Lu�u���_|�������o7����Ba7W�k�U�*���D���֭�L�����$척e�Z�9�S�ݾ���8<���׿�}�}�{'�[r�PB?�k�#P�pLMMm?q��Z���0�R�s3��bk�i��&�-�PM�n�M�X(Q$5�߄���.d��^�}�Dd0��=+��|D�f��D䉞>"T`��ʾ��&if��{V��$�^
������-eMqO<L�"|��@����b��jyRT�J�V9�N�݄�A"�hؚ�H��� �G�7���D������~~)��������ٍ�����[������^�!� �-���h�����L"�4(؃�ԈϦ�o�`������GMo�oz��8p����t�J�]��gsZ����ї^zv[�P�jp�Ģ���d%�6���/	e��Z:�޿?; ��uLLL����?w�ȑ�J-S�{j)͚�M�*�8^~�&�����Z\�ELԫ%S9�fe4$>99��'��i DTW����B�5h�rm, ������x�K�X*:��������ǅ�ԇ��A���h�?��Z�M�b����lJsJ�	���C��X `�T���py�*�v5�Ek��4�wnf�ܰ���������<��+�p��!G.��ƓT,d��zE~�������#!,p�Jж-[���o��nV2_G�l%�u��y(?��ȷ���{;�S+++��+�a�G�V,�Ə��	8�x,��F��d"��E�{��J!��-K%'�L����<�;�
�+�ý�k��fy=c�c�n���o���7��ΛV�My�D�en���;Ѭ}7:�ND�R�|mn ��gq�7�h@�H��B�"� 5ۋ�f���Od�Yɑ!mBqm�qOqT�c߹��IԼ������5���ju�MK�v�h���|ČOiu��:�\��G�X<J��x�4�H$�*MAi���Un���{�j�S��|�\�|���~�����߿/��y���
vb��9��ftt�� ��TO�R��;<`��e�U��P�1��/ܸ�n�M5��v&(���Y��������{߷~�T,�B	H�VIs(U+T���l3�~�8q��<Ĵʽ��&�-{��L<͆Ñt0�;900����z�z�R�|���z�}��<�����h��n���H�J�"h�E%i�H'�Q읪p6g]�Э%s�� 4m�����\���:�T���>h%�h04~�8Pj���	��m#�Ţ@�ᬠ!$�)GK�j��D��.�wB���+��@��P��aK��A������.W�G�B\�\�w��]z����c!HR�h<~��,��E�# �e)��U k4���Y��I���+f��������o���Ͼ޾�ا�pLo�!e���Z���l6������*Ѩ����S�x<���=<8��?��gNOO@?d<*�k^U���$�!JίD�I
	"M��&� �*���m{JS�I���]��F"��d��Ʊ�'�m�𕁁��e�]�9Gp�m� ��SO���C��>h
E����I�!�l�9^��$~�*�.�F���v]ZJs]x[�M�B!_4�����z�Kr\9ٔ�U-s�����'z��3�~�;�1��V.��2NN�[��sXd��>�tg��Npd*O$�̝�ŭ����� _���E:�7��p�y������ ��!�Wj�Wˇ?0##M,�C�����k�O$㔖��܌m}�]����n�u��~�'J��`]��vxvv��b�'�+�+j�J�i{�v��B��V�UmO1���N�e'�<^��3��ypp0��q�#�l��������V���� m�͊�#jOZS�T̒X3�0U�ҁ!u�ŏ��Q���w8$S*b�Ш�9'��=�Z�`p1脲�P0�F'b��ɞD�T��ob��o9��G��B"�+�ܹ��ի��.y�����O�t���l.O�k�#�	���I� ���{ Q�xH�DZKS)����|�Q��G�bl0�'ڮ�1Ec��Zr�TJ��а���~C4:��4�2�J���\��\�]K�N���)�y���D�'�Y�iML��h�R�������c<�J�)}��\;����K�4�[XY���i4I��c��XP�{��$�C��0��R��9�o� _������;.����}ϻf����3���jg%�3��p�T*��lz��K�������`�/��;����
>�78�`(8�;�C��?Gbї�����[�n�W>�����W�����K��8xI�7�M�wV�E���#2��ه��
?R�����c4g���N#��4����6�������U���ێ��^_!t��P��
�pt.	�������M�����山��֭[�����E`yy9��O��裏�?��&�ɑ�=ƩX�ۉ"HkB�VV����w�f��ni�q�)�p|�&���Iknr�5�)$�^�i��s�Y.�<j�uG76�`���+~qw.�h���A֭�Ç�W��U�mX�O����'wD�&.$ ��Vݓ����OD���xR
�&=*qف    IDAT;?O�k�\�0>�6�x�"\(�����Qk>F>s�i��<}��P)�r�X��/��s�|��_ܿ�~?��7���A	�<⿴��&�^�����(vS�M�>��sc��A�:�||P�4W:��){��t_o�B(>�F��CυB�o��$�������,���_���N�<�S�S�/�Z�܃�����.�)�J!X�M.��̇qQp�M�M����ΡL��l�M���6r_O�Q�>+��n!cU ��!	�-ז"H����pg�I���L,�	�G��۹m������={����6Y��^XX��裏:t�p��?n��g�x},��*D���L�	}��IW�:���/c�H�4J���b!!Y|k�R��G؄�� r�QE8���׬�+�hܹ袝����8����q=
���>%�:���r�.'��<q)��I�=v��J�;�3@|�I�T���b���MEB��Z��٣9p�� Y�h��Q�r�\���ٗS�����Pk�f㪫��Ͽ�k����r꠾%��)����l�+S�s���p[C��D;ǰ�Ե�7��"��j�'������a`�b�@ 3��3��I:�S^Ǚ���ϝ81q�W��՟C�ǥ�r�l'��A�k7� ���R��U���1���$��ۆ͟Ь�OAL���������m:g�!�̫�"b�&�*��ng!v\W���#�.�30�G��� ��!����-z<������D<~h��gwm���/�hbǎ��u��mS�������>=���'���D4�,L�$8�wk��4U��TV�����v�o8,V�J��B��C�	�٬��y���=I�>KZ{���na�������w�;&D����p���T-#���N�ז����\���s��V)uL�xMb��a��a�b �:ձg�\V�jۻB�	���>��.�׍��>�t6��M��q+{���ÿ�џ���p:�ׅ����̾	>���ſ��[��S���č�I4m<8�@��H�]$�f�D��	PF)Dމ$v��)�{q�r�
bBIh�h����@�<�X�T��n�I��O�����?�W�?�W5�-S*jc�L��J�D�9�����'i���݂Ƅ(y9�ݫ�R��鐳��a���Q(r����+k�q�R��ﱂ�b5
������{�n��Loooj��=o�@���������ff�C�<�y饗H ��gt���`�+�� /<ߛDZZ��(��K���@� 6٧�����֍-@�D�i}�W��0V}�R���-�:=h�VX��{��Q4}!q񍋫@���e6[��9���R b�
wh�b۩��u.�	�C�w�
hr��*����M��q��O�;� `1Hy�6�i5j�=����v�TN��������@�����C���_~�������g��ӫ�m���6�����l����˟�VS%L]�d��1�/:\��J�H��9E�֑�S���q�����!���7w��4��u���$)>E�����;�)Ixh�lt� L�^�y��6"Y �ȁ��Ϸ�l�QK-o1�c��N%-��e)�L�A�� #���O�4�t�b>�=��dx$���Y��4E�u`���cIJB3�>�ׄC��x,>�ӗ|eӦч�]���mc�]|���4+�\n幹��g�y��bj9q��Is��!�'^(W��-�m����S!��Q�����K��
	K���A�X�� �7�A{����?-1�Cګ"����@��)�FõB�Xd?I=vH H��^��8.�O�W@��NI��(\Jd����J���h�2�OJaC[T۰c�d`�o��4��Ć�lE9q`.�7�9ܴ���Hq+�&���w�Ѩ�M7�wۏ��n�i�\�'�יA@	�������n�c���R�K@��$-C���6��#�N&b�}�Ӹ$�g��Gׂ�A��^+��]�<�� h*s��pi�y�/��2�B�$=�)Pw)	�$�6H9����M�����p0B���nK`J;ƎCfB1s����87�n|A�Y\Z4�j�@hPЖ1�W�Э?��6ߝb��Ra�(��6��A����� n��P�	ރp3<<Lc�{�6�kqS�|��R��4�:[J�>�]N1��3�L�_x|tx�m�vL^w��]sH...ƞ{�#�K�Q�'~jʼ��+fzn�]=�(r.���'��*�Y��\�M>4�w�@^��MB���Fػ�{ި�
�����-�&hh�$��Z��k����Ĳ#㗨ur�PM��	�X��5"�X� �d�U�j���*G�FpI@8�>���v�@`�<| K���*i��@����2%��zmj,Nx�dl���4>��/�l�g�u��U��^�q��ި�~���X,^������B��ds�add�$e���&
���[�Z�m&|���&�ԛ�g�@qJ�җ%"�r�j���!���g�ΛM#-�E����`4l�ՊY��q���3_*��ߡ��5�t�y�>zU��<*�5a�9��@�Mt��T�z�Z`���\Bа8P^�#��5�hCp�n^Mr����5�f���ӧ����8�y�64pцD�B42L��7,!�X��~0^�R�!���E�q��ǚJD�����������q߮�??::p�����N�RW.g�&�Y���'N�0K��MQQ1ህ{)�+�u��A���aN"��]�E���,	(l!�dm$n
��+,)�*����F�=
�t	�b�k���4f������:^b��%�{������{s�CJ�BC��ꔻu���Ƽ�%r\�8��������
&{�!���؂�X� � 7��=��1�e��a�>O��W�u����Ky��C��F@	���.���iqq�'OO��Rȓf
�5L`×�o�G�w������]~���:2OV�T��S��'��Q�
(��M����G�`7�i��_��A;���5}=�fv~��x���7��e���M��j��J�8��A_g��q�[u��$2f9��D�+��̋MHmJW��K��B�3�.��� �xa����+�W�@�|�(Y:8�O��ѣG;�M�_�Ұ ��w�ttt��%���8б {��|�����B8<��Nm|l���g���Nn۶i�>���O��ɉ�9��@MP
�"�'V
\:4�����hq�f0�5�! I��4�O�b�UY��j73�]wǆt���'�kb�@��E��<(�b���mIVl'b!�G��!��ǘX$J��|�t�M(�u�1.Q����!~n��T�c�>��G{U����`&М�	4�Ņ9"~���J�P��A��b������ـkᚸ?�Hp�7r�����H�<��w���?�����٥������-��=77�o�͐V\�ӗd�q�F���۩U�/"G����
��<�t0H����^��[=<���EXc���7�?����[��@�efⴗj�+��0��`���dT���R:e�l�B�M��D�c8�@t8LN����0o�|��an��̵6/X~����G|� t���H�v��Y��5�]�@d����y�w$7##�&�ҳ�:;�)1>T�_��8�N����fi�X�I����p���\�6|ד�� htкD���|�H,<7�a��Ʊ����o���b1gr=j�S'N�x��+OO��$0W�X@D@e��`KP���P�������C�D�ZA��#�5��*#{���s!�7@�G,��@�qb�nX ՑGx���;�Q����	>�%��ɿm��(�
�nv���t��E��"QT?�,i�o!l���{��m���
&�b�,j�J@;���w���Z���%u�',d�$�����Q£Qc�G�x����[?����?�۷O�-�c8[�SB?[Ⱦ�u�fSLOO�?u�z��&���A载=�m�rh�WM�,}��V뵾b���~4��j25��383��s���y���1�OL&<?k�T��3������V#?�
s�&>�x@�߼�̏8�@�8����Cd��pv[�y�#�����(b"xK�yo�<�SnBGP]:�Dc���0�
��f��f||�1��YY�vL�X\8�?T�9���~u����He5+�i#����>y����~ᇂ��E"���$�5�4��Z�FF7<��-�pݵW}uϞ=�s�m_�v?��M���EA� ~�\�\��hQ�#K)r�h�����`1G�� �-����{�D&�vL��s	�s	��\8d����-�s������?�]ΤP�-)�����5%a-�3Ǐ5�R���S�`�����¬V���6�{O/}?!��
�p�[�~0������xh�~_�L�� �:[�{� Ev}OĦ��������+_[/�H�qfPB?38��LM�=699y-�E$�y�f���qn۸�k5t�ݭ�Pz�{���>�:����4\���d�%��_��y���[�]iz9/��"�8���=8����"�	Z/\pZ8`�bS�Z���������č 4��'��?`�>�no6��Q����I"�Gy�8d���J:����A+��$�ym�0B���7H��%;qxB`)`�:?l�3����"��kA(���6� � ��!�C�k�	~~�CCC��|�-�����C�{ӝ�7NLL��|���&��xb(�:���r&��P�y^�1C��:K e��Z��1yN��ˎ�Ʀ�aO{�A;ȗ��i޶ҡ�: ��a��~q&q.A,�օ��?;�#Ƒ]N���3?3K�J)F�'MO��s�T\_�1�v:G����:2D�ľ�Hx�w���r��~�@΄Ns�X�;�A�b�h�4A��Q�>h��	��h���7��g��\����������9F��驇O�:����	�?C��CC�I��i�����砟UɜU9��5�t�T�*`�|gfS���.s��	j���]t���^��o��&H��/�D�$ƍ	��B�H�#>��I���A%ZX���)]���f��&֎%`���`��1��a��3W��̌��:M&��0j��}	�R���L�c�������˹7���6�k��aӦMT���ą����Dǚ�X�P�u�!-�pC�,�� �l��I�\�f1���$a\�@X������w��������{��ѷ���K���LrC�"i�7��+Ȧ��1�B��a��6�m����=����檖��xH�c�r�w���?���S�2�2�ʾ_6ڑb���� 7����M�X�}s<������n� �@Pq��������SXG�+"r����)�T곋uG�$�c!s���=�����`7�����I ��#�.������'~�O���z�֜�1(��\_�OO~��ɉ�<v�i{B� �H�U�@��kB_�ǁD�]��������]�)��{�y��;��33;���6/W���õ�Q�M4����%n�-��Д�g��q�H�>r�b����'�SZ��r����#�j���gN�E ���W��ԔYX�#�ɲN��+�r�)V��ͱcG(/�$|��7��0N�; �P��ݻ�k`ךD�>ֳP�&�r۶m��`�k�N��ad#W���f|���u.���S�3�h�����c����������?��v���w?���Ͼmvf�0@� 	�$_���eE`��D򲉴m�!��Qs��Z����e��5q#Y_��wR���8�α`��� OǇ�.͊��^��>M��)0������	��
R�@m��'�C3���&�����Ёe���"��0#{n���P\���3��\8lF�7<r��}?���|��y�&z�s���9 �}���������֑#G(h��h���߈Dt�إf�ZmQ�E�x^�����!B��c��/���P�,� `�4���#�9�����{���=_x�t �'`mׅ���Ϡ|s�?E付VE�p��V'�� $� m�
,~V}�x����&��`R�S.�;��M�{�n32<F�r ���������[�n%d��P����X�뮻��kM�j�ҽ�c�`.��N����<Yd@�r0����Ü|����K����B��l68H�����{>�K?���xwn���b���/�:r����}��;fg�)�#:��)��O���H�%
��$���ŝ˓X6܂��%k!t�7�߭F�!C���n���s��|vyHM�r�+��N���;�!�[��(����/�j�zh��=a�>m|p?�q~�];d� ��A��D���� ��|�9��s�}���|X���0,H��͛��]7����[~��%���J��o333�މ��_9|�0:�iB���T|A��+�h	�[;\11�9�i�M�D�.�[�e�W�~�y��СEy�ͶM��C)f8,D��/O̅��rA�z]z�t�n.�h^��@�bJ��C��
��w�n�CP	��\z:�<�CFJ�ͅsJ���Ӥ�#:Zr01oy�[��S>��¬YZbS:f�i.��bʭ��p�B��1�CT�Ν;�Э6(�d��{�o!7
H�?���q�����8AT��4B�>Z\>s:ЩPM��=��.��c��m���s��_;W[]�ffw��ʡ����8�|���\.�)CbM3ւ���|�ȩ�z�d6��� ƁpR�\���zd��ǡ!˾f�՝�|�FiX�c(��-���AZ#�)����9ZsԀ��K� t��A ¨7���xE�o�����8r}�����"��~��Q�&n���H>_=�x��-$ ��Ʒid��+�~����/�¡s�?�>�%�s��T��S��;|��>]�\�&w��y�����BZ�5A��L�h8����G��U��{�u�y��g;�,PY�^�;>g:�Q�Ś�TU���&�t#@���A��Bq���Aadx���qMzr��Y�_W��-)L-��|t�lC
m� D- +%3;=M~�R�	�j;v젒���S�V��`8\�
�����W��/��"�� �B�DD ����8xA��N�Z&<�^?>�F�ܞ=WQ�r�!���V����@C�u�<�Y2���}��o=[[��G^읛�?=;y�����S�����h�\�Ӛؽ����Gf^�w\�� )��ȵ��%����`YY�@��1/i��\^dP�kr��͞Șҹ8 α쨙 >l����^F`$U��)�����C�ۧ���z�*��CA�ЩG���IQ���~��g}��,D����j'��AWޏ��'�y�~��7[����zz�/޵�W]u��n��7u����X��UB?ǫ�n��C�^9x�豫Q�1���!��j�Гd�]�p[C�B�n��k���'���)�������'�"-�jm��*|�6lB�鞵u�l�ϷU�V���C�͌8�qpC��pȂ䓉z#�L���IQ����T��UZϓ���ϥ�+߉�B�N�� �j�B�F�	��}�խ���Ej���Ud׮]d�ŵ@��.���2`���"YZ@d�E�R(D�
��W�0������i�Fs�e�S:��ߺ%t.PX��C@���&��y�{�������ǧ��Rs[�fR�.�/^ZN_��fǫ��H�\��F�E���mt8�-?
�؄^�h��R���]s d�")� ���1�#�j��%����S w
ƀ=)n&�g$�:X/�бs�$`Q�u��Y����@��� T�qЦ籞����`��3��b}����ɑ�g���z�6������mZa�.�4@B��g�i��1Tҙ��[�{,kn����]{�o�~��?��Ͽ1PB?�655����O~�ڹ��N�2�q ��Y��m��U]�rk�w9%0MH�����=��ڰ�E%Vm��D�HC��    IDAT�.�"�	�0ʝ����YSj��C���(�K���i����n�M�g�TcBgS%�c}�����=d�y1�:��177[ҫp(���~~�a�p?��4C�j.�qA�t��x�A�����8	H�&x��1�?��Ŗ�����+�N����+/���k�?�`�?4t(T.�C�\4�*�,�S�����bqG&��|%��R*��Z�����FB��CU%kA����3� 6F�<ዖ� r;5�W�����D�7L�2��ڱ��N��u>���;��z�u�
v��L�1�K~9Y��,��;!�1�+{A4u҆qO����֢PN����%{�yZ�
!d��Xy��i��}��2���	�:��bO���b1��o����{�U�������8�[�#����bd2��S�&�=y���$>=:�N�a�����`s���~���g����t�ܿy߷�?=�X��A䬩J�:j�w�fGP|����ƈ�9X�����B�35��Z*i�.B�y�oZ<N�����u.�+~�R-�Źy"t�Ս��c���9�ܳ�4��qBXa�\��"��:S�
ux�XL� a�Gjv�}����:Z4|h�T(�6rA���ҷ�;�qD7�!�"��@�"�W!՝;w>>44����o�u�َW���i��j��W*Vz�z�Yok�j�^m�k���Qk���E�t���iOB��p����el�:�JC ��k�P.h�'i�.F���Wk)�Z����[�ӶR^��Tƚ��9"w�S.E~�Иmt2��̐�D�Z����s�G����|O��C�&b���G#&�����E�6�h�} bψ�]�&�6�{�W�D��鎜˜���ӛ��Kzd02!���{��=W���v��5����|�R	�<-����5333;;;;(H�.��������o�&��[��9!�r�f���C�����\b��&t"2�zLڕiRU;9hjD��8�H
w����s�X�к��E���-�v����_H�-��\�$�h�p`b.�J�,/��.�M&{���j\�Jq����7\א�bnǜ�do��\�p	j�p��%���c �㳢�$'>�F36f�;�qĻf�<v�d��N��D��6X�iL�Y3>�3-O�|���m^_����Y뇭�_"���`��$@K�%���(+�w��M�Z�Z���r�"�,e.�K+�=��.�Oč^6k�Lߡ���.dP>�B�dTJj�*�>�Sp�i��Y��xLY��H}`�@_?�0��jy)C������VPϾ҉>g�n�V�En�;yO��L�^4��G�r�:�:D��K.��O�������h���t����*���U9y�䭳������U��8,@�[�2�2��˭%t!M�.e����G�f{�)��w�B0Tf��h
0=sC	������Aہ��A������/���Du��[k�8t�	B��Pd�2��ψ����ck	�[�g��M��9�x_� �*Qj3��3������2i𶘌��q�B�ƽ�:������Cx!R��bN�e��̣Jb���|�-&s�np�Q!11;C3��s\'\HH�O�+�8E��1��5�,0����~)"B�9pT:��!. �|U6�.k�ڳ�H]R&t&y�h�Ӷ2�Us��!�H8�Nm}��� S��<d9*�di-�g�|j�d�L9��𲋇�ks�;�[s��
qJ�GЪdn�hA��H�.�U��/p&�bȩv��C!���G���	7�a���B�ݻ.���o���~�����ٽ^o��~�W�ĉ���|�\._�h4�A��+u�#���tܦx�9���"(�N!7h�/�p�|�o��2k�B��f�wQ/�44D#�<\t�A�nQ�>z[��cV��h~��D�~�̑��:TݦW�[�sc�������nB����n$��=���Q��N@l2�x�9]|�Xh�m74�L�K����\9ca�ރ�^(���u�����or ���c�d�nr;\\䕴�GE�c3x�] aKX��6Ok�P�v� ���n��a>�/i����B/0[�.f�	$ȇ����!�SÄ�s1��.,PeVD�����"h�� ۀ"�ml	��,*�Ri�J/[KL�|Ӵ6U��F0l� ��{�[TQ-���5HJ�H3tHI#�H#]҈tw��1t�0JH��=4�p��������<�^g�g�k�w����>%��&���
��f�)���~f�H()�&�6hf�KI1���Q����Q�m�/V59�O�#��s��?C�¯�$��o���W{CaW�W�����M�����.�&Ɍ��E�����%ǎ�^#S�HI������o�%���{V�[�	8[�����6N��Z<��pm�@7���V���hL(������q�잢Ծ��Ĵ��"U�2;uy�,㣈�a(I���u~����g�]C>	�Ķn��>R=�#�:|y����M�i\QQO��8O�C���K⁜wg@�n�#�]���y�{�M;��5	�k�>���L%*V6.�G����2�q� �|g�4�%}�?o��$*^��U����-�����<�E�u.�Z��k��H!f�	Q��|��jf�_|gH�S9�v�j�Dē�d�:R�9�ڭü1`��g���SK����ާ�?�C������f?m�"[��Y�+s��<��{�yY��	�ۜs�E�a��Im�7v��egig���n4���K��Β�\?����hq�!ཻ���˝7Gm�P��/�f�� �&� ����aS�Dl�;-��������K��W���(�Qmò��y�
ۂ{�Ԉw޹�Шv�M����{c≥8�q�k%^m�^͇1]X���1!
o�<Wcxhb \�_"OAQ�/S) ���������(���������U�>Q�|��vc4��=f�Z�-u��H�[�8�:hx!�����o���IL������V'
 � �E8���<���ƥ祿&%Zf�t�w��տ�6���'���L�o	���Ap�isG�Q�1���y��΂ Ɯ�.�0M*Nr'Zu[���S�K$z��%	��4ɀ���F���|�H^}�mc Ǔ���UKt�[N5PM��2��Es����>�&��ˑ��,s��lp�ɡ��m���}�Rl*��"���*�*���~l�J"Q�2`����N��� �8<|-Ί�!���#J*rQ�11]���VZ\抌-��_3J�~��Pi�c�.k�˺1N�]v���./��2�a&#�͡�q�F<Y*IB�I#�v�&�3{�2���C#�C1+�6��0��m�������S��h�o�O#<�z9g��AS���>�n�����h4AU�r���]H��f�
`Il�PY|��4Q^d�x�U�N�����$<A��z��;2M�_j��S�n�4c����v��U�I��A`�Y
�L� �0��a�\~!;�BN���E�O����D��'mG��h
�_�t�������DoB�L����٪\�D;�7��@Ds�O�u����N?��y�m��X����DdSd3��9|R�d��r.t��$apU�89�'o�9{��B�v��"+^!	P��H�]%��A�z�,'՚�g�B\�$���&�@�?Q*����hr����/�~��ᾠ�����I�sh<ZI�`	:%9^���c��s�����b�m���|!���:�̎`����� I��!��g�kT��!>�9�����57l�wr�!��+�O�PG[�i�&
0;�҉��C�)c���g��S���D�S2�yN
;��"���}U�V|m��Y���#�꓊�j�'����I$�~��%����0����a��%	��شw��߬�l�~���&���;m�����I_�t�h�$ng�tCD�/��1e$Tr5��;s�#H��ҫ�ܩB�i�,�(S2b���x��Y��������u����VѺ�fj�;��x�%G��6JvH*|l]x�P�^,eN�E.��j�#4A�A�g"u3n�~���&@��޲K6�$!����<�X��/#�U|(cAZ�m\W=lW�z��L{1�h� ]�ܢ�̲�}�ߟ�v�~+ =������~m��&]�u��"Y�o�N7�D�r��g�\������H���I� x������i�nd*휡�q��q���>�C�e�����>�x�K���i�y؞c7��G��ʿ�6f����D��Q�]÷]}���#�N���:k�Hݦ*	����_�.e�ES��vYA��3� 0JH/U�I_s��a��F(�e|�1a���m~V��u�ٙ�9v4!��ZSv.�1��T�K��v��_©��W��2�I{F�	� ��.�t��r
��n�
jAPk�M'������uO'ϝ_�*0�ݣ����E��0d	H*��ߵN�I��`�@���eKC���t����T{���^�X|f���R��5��Kno|7��u��cz\bou˨�� ��(K]���(�0��"�*�Y�²��k���B "eF��v�d�;�x��Mp;��DR�R�{�5���B��Ԑq�j9R�.�K��o��Y�S͆qs8�"��b��5����	D5�p�����:�R����3���C$I����*�s�o%'�;��t�B�v:��c8K�Y�^t��gD�ذ1�!��i�[�8hFX���e1`� f�m���Ԯ�^ܑ��0�[���N#��1�{����=g�x6�H���A�*�F�M��H���*��/D6O�����a����U��m�@CTCq����q�_�*L�;���*X���E�k�[M����wDeJb�J���_J����q�!:�@���籾����6�LP��Ptv��4ZY��(C���~�LdHm�v��O�Dnz�
U1?c�[�!���B�x>�m�6G^�U�#�]���Z�F^�����k��pd�~_#�ԟq�Տ�}kg�:u�4N)��}�D��AT-m��,�N���2��.�����x�i��DDD��	
�%K��E-'$$�e�ۃ��#O�+JZ��+�����jѭ-.�d���z����6��%�R�H!���R�{?7?G����+�ta��n`Kn����sY��RB�����w��L]a���V�MHM��C\��s��GK=�(ؐ�_��#"�=?�������s�\_J���l�;oE���9j|�qsI�g�|��z�����`��ᙳ�%ό|㭑���b >_S��gǶ���$�
�jj�}��Hʌ���ت�G5�
��x!�<@Q6�k߄[�%T��#Ŋݏ�Mv	��߉n��Kx� M;�(;\�O�;�%�R Y�[ĿGBȠG��הE���5����x��FB � �R8�=-�CP^n��oU�W�2�������m/���/�^�T�'�X�X�cݿ!�z�M�w?�Y�w���$*	Z[�	��)n{Z3P�>ŪƊ{fĠ�J{��n��-�`�w ����gGbP>���0���1]�Aiý��lvvv�ttt7�=�W�F��4K���V�	��cOp�Nj�Bׇipq_8qNIK*S��Д�=i5�RD��
|�5��D�jU_#�FZ�B�
�O?ڴ��c��zEY�8[�cy�� sb9��R�KR���c"b�1-�t8�
�ו�p3����y"�O ��3i�EAJ`
� �?>t` ����F�G���i& ��kZXz|`vIt�v ����$}Dw%A��O!>s��<޷p����* �F.������rg~,����˞���?N�d/�b�oR6�b�:,�Aa)e�eN�}|��P{И�i=n�7� =b,�^].ѵ�F��wg�K�QD��h �}�E�uIU�l�"Z��)�d~�]�&iB�E� ��rW���SJ����NR��;ղ���Z��'K����[_���O�YR��fƀ1�!A>A>���S�����A�w�����xM1x̻6���JLWU�<�RX�8H��]�����ι9�+l��{����3�wa�{$��>�֠�p�:�g�0V؁�WE%E����H� �#\��ߜ��/9A1]���+���~��l�$<��f��=Jz P/Q���}?�Ƽ��pi(4��gV�~����x4�L)���oKh�����5�阏
V�<V�F�{���~����q�Ƃ��������/����_7�~1��2$���/�c1�\���Ѵ14��?��f���M��7+�+�2��N>��RG����)�}��&�M���w��q׆Y�������B_yj2��,d]�15�e4��g�4Wv�b�KvNqB� �D�v��Y6\bF�kt��n�ה�jU�__Y�����Hx�@�;�^#���r�H��}A1�&���(�%%���4��Sa@�Y����ބE5N>%O^��z���+U�f����7��:�9����H8�\ }��w_\�tg�U� |��]�]i�%&���S.b�3���)����5_��)_fMg�#�K�%�5�cZ�T�\L�X���eB�H��dz>�}LIk��2X�رٴ!P�8~�X 3"���[�bD2�u� -)$J}�=z��ÿ��+UJW�/ӕo�%�;�1�@!�s��~�����so�.�S���9�{�2�FU�1��������[^�I>K��L��{�*l�xr/̦ް�G�L�VM�����˖4�I�K��V�/8��������n�g���&?��}�A�sG��h�H-��N껎��7��o�u�U��ÎV�r,����F�v�dk��7cS])��8�9�i\�I�@Nq� �$�F�,=#@�c ��4���Q)�n�|���R�_?�B�(BD���7��G C-�5��(��!��g�;^ �����{��22�������f�����u�X'GYM��s5&�Ӟ����΋�<���K�����Z�3�ZM���f�������6WG�;�.Ή��KK�P�ͦ��Eن����}�Q��ǰQ%��}!K�;��0��0�p��}4���b�e��{����}O�v7'o�Ff�jg��e*gʯ?��5'��È��C�@k<�^��!&Z��,��b+&�ѭM3��x��ܓ�>��nWi��gQf5E�`Q���{	8����t_�"Ѝ�x���g��Is����e�o@�ݑ-ov.�d�{���L2��v?v�#{F��������P�}X���8A�.eD��<^o6jI��Zʹ%�ڨV)K�ήŤ�t��r�It���NM��p��J�E���\�8$
��_/����[�(��(�e�?C5���Z�6��G��C�h����M�Y׍M���E�h��Y�a��m�>a�DF���X�񦩥����y��U��4�jա��ga�h��"�:R���$��QnZ�1~r g�XU�T���5JsԎl����8���~q��\������3F��r��s�Z�AU}an�u�cs���	��,@zݯ��f��)s�ۨy#`�]���ۛ)lC�_h���f*K3S�x�B$��f(�I���l��)?�_�vd��f��<P�'wr"�"�X��G�9�$`����/Yg��S�f���������+ P��JAk�r�&�,�I@	9��y�ܶZ�ɑ;�YI�+˓Ij��J�X_45��m�X�L9A���u�t��+�m2��[��%)�=jf�w�4�ء�0ز�8&�QĬvƚ*.A ?j2d۳��	�fޕ#/Q?ۊ��$v����HK\�wy��Q ��v��;�R1�sd��g�ZlԻ}���kg��C���xQ��K%A;�q�d�7^nN;��؊�L~��q*R�H�͂�sK���﫨�#����ba�?�Y&�'���:���`-��7Mt������
Piv�������m�>���c rz�rG�|�t.Gr�{�sr&��[[�(>G�ARH�z�SX�Ŵ��ӣ2>�vo�m�E6�j�/v�%8�"�l��knz�~}~Q�ciXj��z�w�}����栰�TS�]�*ݲ���v�ˡ�Xg��	k����XƇ�I����#j�J �6տ�n|�ʝ0��MQ��.�I���3DC����_���:�����W��R��6N<obt�������ߤ���^���+ՕTuYޕ�ޥ$;ݾ>�N5�����x��n˿�}Ӣ��Єd��1�O�;X[�_�wv��Ҟ��f�S5)�yc}׫�s��;��}�$M���y���X�jc��/̶wk�����a�=�Ì�	�z����a���i����;::322$��L<�bq����c-������<�+"�
�D���dt�UX�F	0C�Q�hڡ66�פ�V��o�NT*��[S��� Vݢ5da]X�L�Is'}}k��=[�$w]v���P�,�gy5T�QU�n�q�޻���d�ʖ�jUITQo�׾t1�@];q��b(��"Z��ǉ���[B_qi�{�t�̇m�������
f/�*к�𴲽ܴ�&�~���|R���{���7���·��0�}h���l4Jt�`Pit=�Y@ ����x��Ը�nS���-b��ֱ��ذ����q-�"˯k�&�Z�`��%A(�UC/�G���D���)}����]Թ�v:W�>�!*ـ7G�!��X�{��ʣÂ{Ȯ�v����j��H!!�����{x���pwC�{����{Ш����^\���yqw*��������n��hz���a��=�nz|�ǟ�E�!�`(��	N��(���ǹ�O��Ҧ(U(��Q����j��δ�:�0:"z�dy(zR��0|�W�e�176���!��[Ŗ�1|������^-���/xb��sвǾ�����,?�Ia�';<"�)���? 8�c����Q�k��1}`�� O,�^�N�6���>2�$���2<�<��i����(�ɔ�����#����<�eZ��`�޵��QW��+ZG�PK   Ԣ�W�@͎� �� /   images/633b3a04-5760-46d4-a0cc-eb31fb771ebb.png��WQ����Npwww������$����C����0�라�9��w��aV�����]�WO���$��D��*+#�
y�� �elq+��tS����$:�� ���U�6<�OU_x�zab���F&������$���]G�v�;�$j)����Ϛ�Ѧ!_� �7������]��~������{BS,g�G�G�>Ao�߈B�������c� �B���'c��1* ��  ����
_�$��'gr���v���	��e(B�O h���� 1�P��L�=���1���&�JDAN��ύ 6N�������?��?1����ˀ���t�Q����y}�2u��ŢB�菷�]�o�᱗2��^>q�cggsl�n��3����--��s#�W8��Q��*�+���)y|"c	��	�/�֎!�U,�ؓ��J��Ջ
�E��D����F���"�uzs�AZd���oU~��ӳ�ʃ�tG޳ځ�tn'C5uul�}7�t���� �+��o�t����_��t�sw�Od������E8U����8~���-��A+|��8�e{.�E˚��v�"K�mǄ��*1���=�b}ʡ���|��ZU_n��z� i��4(Y��<fO&��ʻ��̶�6N��x��l�"I
h�\�F��u|��G�h�U��$��*z��ȼ������".\��A͊J%f�RR�G�D3�1�Y	�����W ?)���w0{�pC
)oK�}�7����,��Jx�'=q�=0G>��~@VI����ͫ~�*�Ϗz���s8�e-"?���\�n�8����Iy���)�s�y��gڭ�֙�h�YZ���7fr� 2bK=�c��x-�k��߉�n�f���QF�����E3ӽ�l�]>����U;�l�n:��|�B��-m��6�P:i����%���<_<k�:
kY>
��qI�|��Ŀ�����o�n[Q��r\o]�й�0�3>>3�����a���������7��8�(�Z���E���or�{A����G�L��ܦ�|��Ć���D���}���c�(S:��W��5HMIy�=���p5-�?�P�����{-ư�
z�����rxV,xB�ٺ�*���h>�N�`C�y �c3��nⶌ���+�>��QE�Һ��"yʔB���&>���)r���/�c����d�[l��dde��m抑WmMLv��2���4��Ao�ojI���.�2�r��Բ5x������/0}q�#Ε3�B6uzj+O/�,v��@Ӻr����0?/:ٚM�O�u士����'懡�00�����f�+�d�`�1�W�b�͸aſ�&9��nm��om;���������z�FŨf�����?���jP�w!k?[��*��E���"�\��c�����m�S��������9��dz8��-�.?�߇?�BI��U�x������8x:��ޘ��!K�3��?�(o�w4�h�;$��$&'��rrz����$�{���7�-�����'s��c�,|bA�����tΛ�������II��Ϊ�>���X��g+*�?(�Ѕ�ߣ�kn�����?q�!I��."D@	�WL�<����Ї�3}M���E]�n7�0��;���r�:�Rt�Y�u��L��^*�y�i8o��~K�p���)��ms;:쾽�)�v\�`!B��TW�g���ךPgŤ�ؾ�+&գQ����}Ul�S ��+��L�t��)>�=�����|=�8=�;�pzu]�����,�� �k���f����M��҂��h9���\H���3a��o�=��1�̝��4*�Pb%(��q�Ӿ������:�� x�=بdj�v�JD&��]G1D��������c�Vy����)w�X|k27�0��SVHY��^���S V��"+�ֳ����ss��&��{1�+���T�!y�7�!���O�1����Y:�^[t8\X22�����"B��΋f�I�ޥ��OE��#�ș\��[Mu�(Z{�D��Bak`G]vJ �s%��b�"�
2~A-<�e&t@��?��@N?t&���g�����q���6.~��9�x^�EY���f����~�a8^��zNt�[UzTȻ�fY��\�����cd8�P�R�i�,���'Fr-��O3))i"@(G�+����9�)�r&�"&�.l��G��=\ˊ=Z���F����d�vo�gs���3�wuf��br�_�w��'Y[4ׇM�׾�$H� 
�G_q��G�ȁ�*Ú��j�%ޝp����
9��p��j�>=[������G�����h\�b[�WX�_? �*dL���:̤jDs��D��Y~;�ԋ[;Y�s��,�Qk),��oh���9���M���9�+Q���YW�o��%?6
�e���%]j�_9Xkvd�F">wmsU�ȸXo�{�PŎI���4��EˇN��{�(��=�`��v�Z�U�xV��U䳴�<WN�V�h���@��xל4���(�?�@T���;���_Ь�[�!���9](��=)�0g����pX߼+mɧ�\�4Ve4�V4׻o%rz�=x�G�ٗXb�8����vd<���q��7=��+E/����$�g��Ic�.ˣ�Mq���H���=�����%p��R򂅅���Ӽp
���O�PB���1<�Z�T�^�Qz����S��DIt����!����?�k=Q������ោO,))!���S�q!���H~yl�XԘsi>��]��i�^RY'�[���=�Pɓ>M�Č�>����+QCʶ�fNAR?�I����'l6��ώ-~�`��>��x�����P3�a���8�9�6��~jv�c�\ZtG�_�M��c������n���5�d��/x�,����X��\q������Ch\�gP��H���j_;qw�WT���~j8����k�V�,m�'أ w��G!�5r��V��iH��Ag�U�1Z�ԯ
�ɕ�g�oUDl[����U�Pͳ��l0 �O�w�q��T���_O�9�ؿ0;�{D���ab_=�re��r�Z8�ת �L������hs��N�|�߁�X��D�>A�-�U��LDhN.��ջDd�Ngŷ|NR�K�Ç���6ۅ򁘘��h	
i���AeQ�rxi��~v�ő�PLVd�J:����*A)�)L�:�9�ZrD�:���Q��p-������777��[�o�������#�TU�`�䀝#�K�|�[7��h��b�J4�U45G(��Ҩ�� ��7���=�3��m%����A���hZ�q�<c�Z�,��ƑR�)hX��+L��|�*�'��"�G���7B
M{[���pÊ�JP�J�
ns�k�5�|D�>>>N��'I����5\]���V..W��2�U#{6���7�() ��g��Y~B4c�I���+)٫�+�_�`d+SHTo��e�8&��P�V{~eyu5�ݓ?ab��ׯ�_��/�Ԕx���)'_瓗�s\o^T�(ͭ��!N��<��ܽ>Z䚖��6U/e�(�v�l�����D_ߞ !��jl�$J�<���2�������iRǊXbȘ�<�џI6�� c�U'A����.���ͼ��O�*��.P�(!�����I�����=qK�Dv��PG����ұ�$=t��5���0���s(h�W��Žp�b��2"�{�]�\�Ai}@�yVH��`#(�D�<���P*rU�8?����~"b��`9q�u<m"z4��"ϻ!��S���\��L^7�ɬ�C����aSK��)��n8da������nܱ~��(��9��n����i�ō�M����H��Y{�]���$o��\
��K��,T��#G��X��/��vOA��.��K���[T^H�
Љq�$�k������p�V����6���M*x	����k#�q5�`/����� ���K "�2(��P��&�)��:2p6&NcO8������э����S�H��b�	��J���῏��
�� ��r9©��T��6�H���ٕ�G��5
�$S#����+�1Kx�|��+�	&�j��B �C7~됂���Z(�,��"��]�m�ף�J�h�H`>l�(fp90Plt�4���"��2\�sP	1��b@���u���?���nn �63��C�'	�Q�-rȕ #In�c��'������� 2��3v�Bx��&�ϩT2��X�w��PhA*`��Xywm~��8����+�D.�]�w��]~^Mx5�]^%�G �ڋ�6�E��ʍ�@5�?��24�a�����[�2���XaĿ2�	��FA���J�����,���k���H��|	1�|jc�X�EPp�Ab��$��:����Wv����'���.Uc����Eh�Qg���ڴ�4�C�{�	.����af�Ϩ�b'6q;�F��vؿ;N��TҊD��f�W>TvH��hMvH/���ᓹ��-��!����K/G�o��o�.f~_PjmI��j��w�=�A�6�sŊV���u�2?��.�h�����ƒU]�@�ɕn�ut;m���菰��
X���x�A1��W�S9�|eF�CS�*�u�A%F�AyT�~���iME�$E5N\zT&�9�)N$䛪�m�{hK��iR��v��?a��s�����CK�'�Q��v�u�-mBһ#4��b����"��Z<�* �!4��o�eӴ��6@btl�H�̢�#`ѫլ��tA�@0��ّ�2�*�ݎ;��"t�qx��bs[�ъ� � sɓ�K���m�X���u��m`'RJʃX� ���ARZ�V=�,�g�{D�b����9K�**+��K� ĪF%�t�K��!SB� ���`� i	��u䑩�7c����Č5sq�X���H�؜\��ɥ��}�,H�1߾��<��[�+�N]�y�c���Y��E�y���h+�	��m��,*�����lW�y��Ѻ��	Z�����7�:^2
rH�@���%jO����K-	u�8�x����1|$��;���'mf3 |��P��'B�%.!����l��Q��v�_�8m������	�ɟ�B��f���c1m���W|HM|-��A&���._��������y�r�#�D���t7�'M�0h_򄟏�A[�VP!�62�P.�}ߏWu�������Xm�=��8S��TK�"�JK����p�=���-,���-ƒ7j]Fߋmt9MM(�{%�����)W�a��#�B������u4ǂ�n�J�UB]��_?j�P���"sJ�#�O���n��OV�VYɒgz����ϧ�{o[ܚ��&M��_���L2d˱EDl�uE�D�hg��04b��e}t����<u��I��7���3��[ŴEC���%�G��v}�#<���t*H��$/0 [�g�]��҂�?;��K�[��FC~�rI�J~#�U��WSe �w��|�y�\7�11Ĩ��Uyac?����h�
����Ę��wT��H<qTH0�Ɔz�'��J��VEv�g��H�~77/7��Q�>�/KP���&'Дkx;��c�Ro��C���,�p���Uh�f
�&vB<����������t��l������&;<\O;ew�oI%���l)�tPS���h���xZ1g���Wi?�CҀ�ī�#�~4'[9
���N�2�-��=27 64�i��!v�;2�ۇ���������\�11N*]]��ɗeݷ>��L%�/�Q0g\~v�������(B�M���XX����mG�2a��K��.w%emڡDD�eE`bd�dW�@1���-U�g�8V��x��"�A����vGJ���V������"�;/w?n�V�.�xeۭeZ���MKlc<;��	]�0����5C��Nk������,���O��H��Be&�[��,�l�U�2b7�nB�������HR)��M��cE���`�A����T�5z{��*��d��d��	�iڪ�*�#�6�"���?���
�RÕ��p����A�.�xS��e�p8���Ft��W���5=�0��_0���SN+�!���v"� ��>�X
J>�	�O���#{���� h���;��T!n`�ԝ7q�VYV�VI^q�D�*�U�� L+���Eh�-�'�����u#
��1C��"d??E�g����������[�l^��,p�UUMDI�f�P��'%��ݜ�W����W�:6	-�T��tjW �r�*$9:�+j\f:,������I�/غ'�>��O�[��Yvh9�r�`�C�Ŏo'���fJl�C�'��[Em=lgF(��x�O�1�r�\�z�v�!.q�y��\=�A�	T�IҺoM>O����%�c6�����:�bXv�dqFA�-3f�O��L8%���yq䱗�i<�A^�6p��2Z#�F:8)����
Ym(t-FӁ��؛�����d����A�1�����8���=��L1��E��B����p��ԇZE��%���EZ��7� �!���
U�x�יK[�S-X�'R.'�K�\P����lJFp ��`"��{r�$��m_b\T������a�"���P�����P�E�j��yC1�Ց�����7��|Z����k��	��x��Z����b�"["��h���etFE�>::�^���=��1F�ttt��C��4P��P����{�礁��1'''�&��m�6��l��R�a����P����+_��m�9F���c��U��{Y��[Ο��2ۋF*u��V�B�e�[#�jF{�!q��w�]�/�����v�h��3����hd��o/�gv������W+:�_���99C��ޞ��n���
�R/��bjvt^Apyv�@�?�5;���_IE�3���\W%6�|��	�ύ��r�h��;
�t���J�Ak[Iod�_眠�%�7Õ)"���щaj?����Q��g)���_��g^1��{�;@�f�C><M����� ��繠ў���2�A���q
O~��ٟ����z3%6���!�k�cx�XU!#p�MYo攅��z��6/Х�>��!�M�C�+v��.�V5B�Fv/	J����\\��#'��S2��5~�63���F
:����o�0a$z�����t�^<�+��00;77GβM`mڪ%)�Bd���'�#�����΃䌑W��ݡ�,prP9o�
\�+fԲ_k���M�8s�m�]�-���xfi�sR"�AĒ@Ą��fƤ�P��q�G���^<L��o�`عLᝉ,�6`Vlf�����ye���xu��;qm�n	z���9����`�������ㄷ�˹�	 SV��s�<��[Uz-�r�}�C������?5�nCVu���Z/V����r�}�O�
\��~�}�4J��F*�Wʱ�rѻ_��ah@��17w�4�Y�{J�!������H����\�T*+hB�̙�蔞&����o��?.D��&	���)k-N-��O`�^����S����[m��-:7�)u3ˍ��1Z8����'vKB��E-��?��ͼ�wvr/��M���%�Y����{,lۍ�>(�Ƀ1����x"�;���  ��NE8"&�Ov��B:���=+ē�k�H�,X����q^���g	=���/C�u����/�STb��M<��Vs뢦��U*���n��)�$��h����"���������F�����������ӁMZh��u��9/��0�1N�J���O�΋]y���w����I�����+���J�Hp��2����A#%%���u�ng 2ȋ�����
Ζ3������f��Rx�n����aKjkk,�%��LuX-ךЃ�:���z[ª}�=J"E<��U�m�I:#	�n�/�W��E��K?8;g��Y
d���b~w�dh���:bJ������H�b%�q#��n����Uxn���������a�d 篗��c������BXG'�F��X�V�V�=���t�ܒ�-n�X�D��c��c�i���E0�"6�~|7`���	K�;A)*,����ٸ��g�Z&e@��${��~.����k)��cuq�r�U��l(�լd�����e��f}Dv{g�H��/�a�EY`�OK��dd�A��
qR���C'y}�!�9=%��X�rz;<pFO�9�e�P��
�w�
Қe������p�h]X�vZ�"/hJ����l�{ߙ'~)g:�Ε��cyVS�Κ���F������Ʃ��s:��ypW5K�l�"d�R�/D��ƺ'ɂt�ulBܱ���%��s�����
�¬#�bWeRE�q�E������}��5���J>�Xf؈�����|���x��e�m���YҰ���L�FH(�Z	�'F-Y��C/�-�=�7�5$?��,;S��FGL���gl�{������qR7j]��{W�Ƃl�ċ�����nUO-7�{��q��\rr�ү�a b4-�s;�F�+W�������/�-�������f����+a���Y8&��z�/��:UӖ�h�'h�����*ǟk��E=Z0e܌�u6���m��\G3;�N`@�Y�$G��x�?q��"~��[&��m�?	zzhhnv"�{����>=ڵ8n��?]�0�y���`�Z�͖�1��� a�</��'�i��B��{ZG�cY�B���P�O��z�ǚM�u	?~����b�>��}�U�L��W*���"�[���[
�y���Y���f�f��D�j�K���"��l�!f����:m7��C�P���7�.p �\�_AI:��7Ի�;���NI�Z�+�%�o�O"���&X���sEF�u��=m[عT�σdm�^�Lڬ��K��瞸�tN���3�e�H�9~�����Z��ox���d���|�Db�<2nk�i�6ZN�},/��n�Q�S�r����dа�=���b��ic�u�y����)���S�j��c³ئX����W�C/�p�����[$�)���� �z&lmZX���Юɭ G���6�/2hz7�ꋹ
`���ť�~)��ya���I��Q=f�O�&�ܮ��.����kx�<�)�JS��/F?�k��,��ԬB���m��F�I�J����Y�p-q�3�-Q���w��A��ͳ�O��^�`�0�gPK��)���l�,ˊK��d� l�YU�٥۶K�70�}��;]�;M�J-.�_�=q�����+����7��=./���팂M�����EI,����n��;V�-�s�e/π�N����j�W�q�j�[��C�;H�a̙G�8�2~$)ݶemóccX���DJ/g�&_�BΝ�_�	)���/�7W����AD#��6�G�6��
����#�x_�;WՙW jV��oN�\�Q��%_jdXSZZZM�ۤ��� ���9ɥ�x&o�vW˖��MrU���)ȳ��5'�
����\��y? ��|���ϰ+�"���9�!:��^f����n�}��\�ڿ�j*� ����_�/���O�+��z#�V���J�(Ҍz�Hbj��q������!�R(c5�IA������,p�Pp�ؾ����%F�h�A�m��3S�(6��U�C���[��E��YXX�%�ZM
܌s�WTt�%3��ǔ�_�&(���ƛV�N�|ZFl6�D=��YmK���l4&�K�S��~��f�2� �6�[T��B�	v̙�)��H7�e 7j&�К;��a$�z���VF/����5�a�͗������jx�=���������b����.��.W���T�j��˶����T�^/ia�-W,�:��o�$�?m�}��|'V(D�+�`��%~��C�����f�q�ж�ӧ�ŗD�zE�)�����g�8����K�7�V��r��Q���z��y_�Ɍ�-��\Q����O��C�:�GmՓ�T�y�M�qX|��<?�k'c�K�~��#@��Qz�@�u�<����jq8�����qD��-Z?�#ժ�Dml��m��c�!�
;ް��&s�t5I�e�>~ C����\�"�dz8���e]��0�����ܘ�೽Q����b~����r�xj|\�ƹM�����ȩ�nQ���1���l��x�CC���A[+f��U�t����\TOz�/\�8w��l�3�� ��	ƕϴ���W	o�*���Ձ�ͭ/v�q��$?==�P)e+J����!��}��yS��>'S��>�_k������EG�Ɂ����;?�?f{�zQZYc��Ĭ��'�s����|�"��0��z-�i7�5	!�S���X������uӫuֻ+��w��Q{D?�a �e�̟�H[�&��{�6��/��Sl\�\��=c�&	8^��l2��B����̵���ħ�����X�ArU�l9(%hb���-:C��@��Ұbb�����Ob6,�2h ]؞��|�$�����ύ�N���1:95mk�¾e�\�2q�����U2jv��E�=U}}�����\��jv555yn�uo��I5�9�Uˆ�'�ȉ�u�:�J��f�-��`��Pd���/��ga��9B]�m�28�E\D��x��/lmG�B��/5��+����e3���6&���S]�Q��\���sHrB)��)
�
���XI���`��z��t�AEL���M[B���ۈpi���WhɎ������	�g$�^��_�o�[/����>�BllM��l;݆<��⼴���q���[�����{��$s�	����U]� ���bG���x2�+�8dL􆣑�ׯ�)�ȸ�6��V9� �� �z�)n���<<llm(�ù�*��|�FH�B��������Ԛe�iǖ���"�tm�:���&4M�(&5�@U��8{���f�qw��ty�~]e���b��������; ���/vH�&��.�^q=�����]-�I?z��2��k���
/`�T�	�����0�lU���)���3c� ve��� :�@5p����тf���_6j/+0:n�2q����`�����i�!#H:��Nعs�Mb��5�$����Tk�=a��_}�z�:#ʖ^Ӱ��^2l��2#L��>���촇�AI���y��*wܐ��d�p�un+r����h2(�nA���i(�d<[�0��m��ϟ�eeeh�X�q.���r�ڤ�{���Ĝ�^�I �+�C��A�g����`U;v��<��,%#����#O`�JA�<����D�8���0�kv]��QS�Y,S6I%�:HR�����ؽv��~|���e{{<#V�'��j.2W�\�� 4&w��d\T�H.h�����ܶP��A����:���'Vpy@�rnWܘ��+�rw:ם:A�s�32w�Z��5�Ȑ*���ٹ`��B�R���X�f5|Y�.�jN����mUy9�
�ჟZ��ۡ/K���݇rC�c������{�<���I��S�4��6�I�A�.)�c�܇&�}6��i*�KW���n$������a�:DD-yk���4c�������Y*��f&��M?Ǣ9�6��	=�;A����l0�Vl���]�����-j(T��l�ahB.�OXh�Uq��bZ�I\oڹ�n}�@���ou��U�0V�;�;���ժҁW�?
Q�$)-mG������&�[�9D���+(���l�=Ec��vGd�!~�'%���=y���\A���ߴ!��VE/I��x�:_T��_	�l�L~ԋ�J�.�0�Q��4k��zx(j.�K��n�bq�J9�?�R�����9B˫	�d����E��xX2���v��9e�u͡�S7���)��p�\N�	`F�Ñ�:�
���Ïș�?BJ�������A�#����#��<�|2�@$D���洌/k���B�-d���C�{�y?2ty��k��Z�%7��$S��v�I�^w41�w��H�r:�G{�CT�����;�6����y��mj'�j:Z�Z���@�+��5#��cڞݮG!.�e6�ǀ?��M#\QL+c��>ga��=�Ƃ��Rn=�â����o���S����L#̺s�#o��bĬs�7�牲>�[�C����,����m�Y0��I�"��������Z����ԞG\1w�Ζ��x���o(ι{���\��"甯�)Z�ݦ���$�z�gR�"�u~�.����h��[��v�fqZ,ךd�k����9�M�y_�Ƽ�]Ԕ����`�}GD����pWr�Y����hZC܀�_�8�4�����r���ɶ��2Er��`\��r����?|*��{�mht��ZOV/�y�j�#3��A������F�l;�ͲMIKL�1���t���y4Qzǭp~�w㏄՞�ToAX�=-�)I���K'����?�yW�.��q��0���cV����%P��ʂ ���p��5d�-)*���+�@u�����2��es\o�_���Y��F�x�������3+�Ыq��O�
!V�H�q��˵!@�mq|[��	:]q��~n��O��k��K^��ە�Q���l�ܿ�鴸���X�M��#�A��,��F�(O��tڇ��wz����o��~��b�<]����6�4m��j?��+��+������P8lt�J�*3����ON��Z�;�OKʁ��`zl��hok�����e=T99��]r4�������P�>�C6.=T�	=��5�+\�'��ϣ+����E��;�(�E��{Z
&��xa_�s�Z����@h���}���"��u�;�<{��+h}�P��61trݫ�[.^�ŕ��x�(�g�y�uf� �h���iʄ����2v#t8螽Щ��<���d����n�?A`jjI>[�8ڨЪ�^�lh3���~=q�9)C��D4�C�<NG����#IJ-�ҷa��C��o�ׇ���˕�-�ƘV��ҋ�۹\;�O��¬�?3� �RĚ�զ¬��7��Λ�X�H5$��+@�@��z�^�-��c�Eek��RyB	��Yک�\qO�����B������uw/N�H��u[��^�z�^�(T�`f��Ƃ��>��昮�i8�D#�O/)#4��L^^p�Zn�{,5�g����ݟVj';��gA0���b�g���φ|׮�8�,�A�YzY�H1�'�b�-e��}p�.��K8s%�+���4F�UU �8ܙ�Zt�,$���#=�������V3�PHOe<L2�t�p�h(�k�P&��49���F�ћ׬R;��UM;ct�G���@�Ɩ��Rۥ�ޝ�tltt�7b:�W�,dԑ���Z�]ɚ�VVZ�гC�8�����Uk�/�r�)I����������V��r�Z*3==?��/&)tE�%;��I%�k /|�.<ʰ�pj�(<��6�Nȉ�;�C�א�vaw� 2��)r��42�[�wS�Ѵ�&�����Q��&ҷ�{�v+����)��6�#�/f(��3P����pi�h%�{���5ؚU�h3Ә��ݣnZ�?23z� �Y�xR	$c�!Вj��ԑ�� k�j�$�a�E_GG1K���İ�ZESC��~ew*'�~�r�u�Ґ���5gg��UG�{pE�g �We�j'"�L܈�\ *3�_�b"��h$���g�+�@%�߳��-!H�����G��*WqQa��L�����f���J�j��VVR��ƿ�.��@�/���c�FWW#7��|md��0�!�x<N�I�|{����<�A��>�Ǆ��i�P����/
����w����_��yq\۟����Z��ڎ���_��6o�mX��_��Fr�UU��-T����D��U��]	��mg���z?9�!1#=�Y�a������J֯�:���ЂA)%p#x�`�&����_h[��� ��G�g��yf�J]J!H�L�0�� �i�����+��pt��h�t��466�KZ�ۉ�O�;���e启0Hz��b�B(,j�E�X�艝�|�^��ex��2�DGCs�O�����|��_�T��Ј�wBas��c���ѵ��Q����B�g�g�s�bË��4��9��6��#(b���,�:D[`"L\e6�2@pzl����G��6Ls����D�(pa!�ߝm�|0�5�����m=x��	��~��3����N��|�5dڷo�������y�ƅ<�*hb��J�Bs*�}VV��|]����%�WT"����
YH�8��ܢ�OU�����4d�TCG�	��*3p�aJ�c��e�Rg�(V�l$�Թ7<��"_��k�g��9�^〵�b{C�<��|t>�K��ó�:73>==mY���o֙��H���#3w�r��z��|�����q�2�J�����~��τ��@
��4Y�%�G��Y@Ck{�Fe������Q�l��RPy�
^+�Ҹٞ0����X"��{�	�,_wl��j�@G����|C%���9R��:���0���#l���,U1@����
ef<�uƚ�c�H� �2��w��L%"	�Ms'��/�X��ofyA�Rr��0��IB�������D����"H�J_�
()ߺkz��I�n�Ք���W"�^�:����qP���Ff�2@Q�<��Eڶ��G �
@���Қ-�,�7p,TQ�Yl5�X���< �GV���W��V��#`l��]�'Q:��s�[t�I��)�]���b���A������|��xsYvF�B�[��Ç_�"T�)Y�h ,v�9~�v��4����"%Y�5(���� ���Cv���A&sx Z/4�����}��]�/�C�c�3��^�@��.�f�a��>��o/���@��9���I�{8�����YF�	UAy���IIIeÀ��"��WypF{LX;�I����-//�kjj�Ԕ��AӢ�z�H[�����=��D�cQ+,[!�e8��	����,W���(�;�����G��P٦ܮ��e�+� ��!����;qm��}b���_|�\wc�}�;H�Y�{Ʈ*+k%n����a����W_[N�O��F�g{�e%F �e��Î"��1%bpG}^]�����ȧV)R���b����i\�y���$Ʌ����K�)яܼ��V�a*�8�&��W����#����+�d��a9��$��[W0����l��P��y �\�|���K49��N�h�nu`���b)�@�R��������Ru:�I~A��!��!��8"?�|�q��2�G�#�V�]���r����Q�6;��Ca�ϑ>��I�u�\���I�T2�&6������/���X�d#f..��B¾r0���{�o�-�m�d,�bٕ;<�qx�И=�����W�����6�`����Zpk��q'm6�I��L��ߑ�}$�x�a&_�W��q�|fά������Y.Q>�>�y��.�+�,�ے,�W[3�66.��cv�[e�8'��ȓY�f��&��D�`������fo8Ώ�}�wЋB�֏������ ��ٲI�tr-���j_^��:Wj_�-;��leԶ�_�G�~G���m�J����`���gS�V- !O9����f�� �������4.���oR���-�V�����^�+��	�{�w+؉����Zq�J�8@��0._�G�Na����%SOtI�:S�0�n�{.��R�)˃�������j�Hd���dq���Ǖ�G���=;���c&�ΕQ�R;��qWQӝ�ۓ�d�vB�Y��@pϽ��f���kbe�*v���ֆ�"s��։�0\\�ūX���;��d��	\y��%��u�(��ۓ	�T���,�1@z��O8؞�e�^��,M���)����������@����z�Eq���٢� �3ϗC���x����Sa����^���I~{���i����D�=������K�=�f�--� hY�HIwm���^ʆb���~�U�+_A/��S`�k��'l�{9�P[2-�e�T�7�y�agɈ�z�;!ڢ}�Ɏg�ߕ�L���N﹭���sPpyfy�'�g��T���AZ��P>�������6��HNo������Bs���N�9k�9���NB\{�� �n2(<҇g�ҽ=TK�'!d�6X�C��6����(�����u�.f�?�'��L]������EϚ��tOMM-hJ]Ē�%��1|��N�J�:
	87ܭ<�jh���WH�$=�͑kk1C�mtLT>kY�s����������(�2��&����"�@M��ۯ�������̂
�{STG&�f��˙���$��.A����1��h3�[��Ӣ�m\ń��_��*L���w�M�I�)�&��Z E���X��fn}�l�/���U���l��|��@VYL~ڦ�����>�	��$�K��!�M�i�.xh���2�ͦ[ø-�(�-�R��ŝ��w/���b���!X�p·����<3Ϟ{_��ޓ�:&�4�6#�ޞ���Kt$�$FݽdU�"�O����&|��.[�Q7�e����p��>��ψ����=�-*��!"&�g��ȏ�X�1'<���S̢<��K��C��Դ'���p,� K�4�G���o���
��@.ל���Y�S�T;���k��Qė�l�(��<Z��k��%���	�w!2\�gy0���%9R�Ρs��{�W�����;[CB����g5TT�:xl9ͫi�����6��NUJfe ���=�Y�51(�-m��v�4���Fh��./�F��bȬ�sm]�A�fȱ4��f�ulX��d�`&nS��Z�G��H�;�TӖI��C����)�_�8tp�z���X��4�4O�7�H�skg�j��|�K_[����"�����>�i�M���s= �k�:�X(��pkt��v.�����X�;��QF��(`$q�x�r�8�B��E��1�4��/:�(����L}!�ɽ�����D���>,�ƹib,h�bK��˥NDB2N!�!���=FlYFw!O d�	'��*����|��u�����i��'��:RQ�ժ-,������R����{�_ݛ���\Id��H�C��y8!b_3-���)��+<��{ߵM��m�&0�����矗�]�U~e��zK.6RR>�v]�v�ѿ�b�tRȺBT�"�R�^�AY��x�F�|~�>ѓ,��pQ��M��g	yJ�gɏ�]�Tl���z)f7��sxϣ������&�-2��)u�ʐ�''����u�1�;�X�9g�N܈��ҵ3K���O�m��u��W�:�ށ��\ܾ1�s��rez� !dAlf���T�͡s?K���o�0� H���N�������8[@^�ҽ_���EBO�0������z}�k��!���-������S':�LG�"�'�M�.xw��Y�G%��EJ��)��6˭�AX���|���}���d��F��<,BY/W5��]���F��U� ,�8m��rRL[�?��{7.z�C%l�j�f����d�b��N�\ �6	�m�2+��:�(��7ڸlw|��)A��l�#�'�v�롍����Y�'�Cɑ�韹�VE�\^�h���A��ԕ���rJ��4�RrVVg�\�� �\B��Yφp�r:�^��6]A�F,&��\�ݑ����N�aIw˝�r����*K�ۻ�z鵔}f.�la>o���}<D�bW��*r���lI��I�L����;��N(\QBd7�E��4�(��ׁɖKT�l_�� F���:XϷ�n]��c�X����Y��ͬ-tR�V!��XNF�������V���/|��C�3Ҧ��oV��^cQ2��a˧0��tz_����Ľ|����7��Va�BTsv �q�g���Jc.r��IF*<���<X�K0���.z�.D�<�7T���P2���u�%�B��(�܂�}��ʧÅ~�]9^��3	�9�m�b᏿�m��������*b��;]{��&,�O�K�����Y&�&r�c�`�bK�3�uG"G����Z~s<�������0��e06��V	��m;7Q�Cj�J5 �z�]�Z��*SDx��Vd��`����4���:�Ƴ���k�����t�l\�v"ϫ+?�|{�Ȫ�;;�^�x�Z�8��)�a�����&��yQV:c��Y����ԑ��pLqԐm�;;YT�Ew|��~���%�u��tQ���"�#���G�=�����K�c��l��15$�j�P\7v͋��M�:���g�����M�c*?Jþ�ى#��$Z�����j��t�׳q+Đ���w�&�񜓑��"��xxyA�u�~����Sh�Ol�O2c��~�H�7��#�}� d�\��\���n��ey�#2j',x�-~!����XP��9!�����(a;�w�𾃐�`��풘�a�_����bUT��k3�����9[�'�J��&yd����#�����a
bl�"��8~�\m��#''�w9V7��ן��w�+%�S��Z�#f.��.���D��B����6N�+�;�_��C5�=�R�����O�� ���$�k'��-|b����K�֧��I����֬};d�U�Io��,7���@[;|��$U�1��|H�aA�/���f�����0�����W�����P ��4J��� e��o����\�ݪ���
W�98k��/sQ����F����5_^^FxK�=���� �R<1�����Ut��Fy]퍩we8E�ɘ����C!~�'\�[�����X3bc��!ԫ�͜�D��5�6�|���}�rg���$>���TN��j�M����J��Yw��tS'F��`*K܋�D�Bg�		=x��c'��P!�g̮)�������-�9������y_��Ybbb$�Z^�:�W����F�ӛ"��?D�� �Crʂ���[���41�s�5�U0��K�=����������.���B-��o�P��� ��%��� ��кo�ρ%O����̹��?����)q�'!��w��+ײK6���T������`9e�&��(1@�C3����h����B�^��3|2�����q������xdd$P�Hk��sP�;Y��ߝ���m�w\E+����{�S��?�L,���>]_�|*�D�B<1��5��Ԟ����E����.��p����_o�	�^~y\��d��<6J3k�d�sɜ-���q+���Z87�����G�;P����1aP1��b��C�nڌ�/wc�No5mR8�IS���������^��[ى��Z�ɜ8%6�+��hb�:�s��*��wb����+��:�X͔�����#���D~�_� ��(u���ƕ�R��Eiem��MZυJ��0�h�ސ�k8�Hjhiye�5�Q��v�0!U]w	hKX��Hf
� AKU�;��o�ry���� c�zxt��>p;W��)�_�e��P���DV�Bɻ�@N����'�C����w���/ȴ�]?����h�X�v��#���?n�)�a�͎�hʠ�~��1!;��}\?tF��鵹fzO}c��7<qm;tj�SL��{�����g+Z�awo�Ci�ͽ���ov�Oum{vsm[���������i�&}z�7��U��m���Bz���4�q�Sh�㿘.i�k�,��3%��׏���ht�؟W��XL�Q�1l�=)��Y?s�W��'z�k��^����s�n���9��q�
+�X����>'''}�^�O�Ԏ�
^����i%#5ْ�q2c�ll��M��1�hH:pXZ��>�C�ċ�$�V������KKYp�'fr���=1�f�5�jz�f~f��;�zg`��0iq/eUbc�F�ȴWW_��Uu>��*&"%���Ƭ�{W���F��)m�$���y2��q�
�&r_WRF~��P_C��T�D�(<N�$���i8uc��霨V��g�m�<;t�o}ҷ*s�@{�ƕ�^ں�T���h5qm����tD�(�$_�oÏ�փ����3_s��`�Ln�H+(L��.۾���3�}懞��Y�v#�d�����)�nb�@�"7�z�{N�j�9��u�52_�I,��ܗT���e:U�������2��Z�q�z��ۼ��=ˎ�W��J���1U�U��?��� ������n$�@�W�G�1�N�R��_Af	��د��,�g�G`PCS�<��}aWپ����1���B~��6 ��ǎ�Gu�V�C���C���U��D_��h����g�.Y&�]1���l Ϡ3A����d�����R�Ĉ�D�ʲ��r*2J,�VT٪��1݋��Y�G��2�S���B�	���¦/�	�p�j9�K���t%$e7�����sU,�W�S�5W��S�ˍ-����5	��7�k�fuZ�<s�L>���Aڷ7�]����DKqII�y�#I Qד�ך�p�wp�K������?���E�������Ys���W9I[��^�x��w���`�ڪp?�Y�/JӺEH;���L�*�E��:	s����9fi{�ϏP���������a�y�o:*��.�Y�hi�Jr��y��m�쁖:h83&��������:�F�զI_�z�[8N����䍋��`,�e������M`�IIK�HK��x��z�̾��v	T����0�q9'fU���cX��2��zPm��&6=��,�,�2�)�������ϭ��$D�9A�������p���� lBVTd�9�V��.����+ɣ7�ڵ���Ç!�qc
�_B�3�:k��)�(:հ���qM��P�8�l�� ��nUɻN>��uuh�A��F�����'&�EϚ��Y��/#GvE4br
��%�X��l��G�]�x>���Z�5VYi&�a�(1����$�VҤ�)q�5�TbS�6�JKO<���tz��vN�I�/�V�Fd����O$~��u�e��V��=CI��WW"�k��	�gm�pA�ۆ>�A��Pr���͵p��XD�z����N0��D�}yi>eX�Vh�7Hp�� ����%Y����v�j�
ՑG΂*�{�\�Ys�[4���>I!����5�7⢒ԕ��Mȳ;5�ң~QW�&F��	^g��[8@�)JM@@}������t��GՁ#kl�r���nʑ"��Z�3�y��{���ƕr��8@�
��ָx�\942�#�̑��Ѓٟ��2E,[)��@� �.<<|��ٷ�b����t�����Ӥ�f� �ƃ�"��|�*i�ûꖆ�%�*`�{^b�J��o��O�U(Bj* ����4�c����s��C�@%��̦X`�<���2�>l��Zڥ�.R���/�۾�j����=%��L˴=L�q������˛%zrVޒ���1��a���#���D���"΄"��k�bu4~��N�2麃lCE�s�U[�����78����[n���GJ?��pyDz��<_��~m��9��R'li�{b���` ۉ�>{�����ʈ�2��x �q����������Z�(cV�s'M����&\u�$����>(|~W��W�x7!�Y�6�2�u~˸+�&;��F+��F���w���aP٠ �e��_�"�MMMeW�䪾��W�FK;!|erf��';��pڡh�I��6����>c��cޢ������#��b釮n$@��˰k���()���Ҿ�f9�YҖO(,���q�ESF6F���B���tZy?������-�g�4�Uut��Ŝ�[��r�g
/|�+�J���C�~��ՑS�kS+��#����s^�ó�KN�_�/�����3�v��2�}����х�::�:���o�M~\C&�_]��Ḭ,K*���$��'�~���>�]G������{�����#&�m�t�8!���e�]nO*O�?���.���W"*e[d�R�A�E߻T��� nUUxI���F�kp��:+oQ��+�q��(���l���q�[��#c����Эw��K#��5�kS��h
�,ܳ(^	�ֿǳ:���Ӥ�-��cW�8�w!��q��r�d�O��:��HeO,1-��k��:��r�Dv#��p
����٪�.�s���c���dQg�wǙ/�%9L�,��]�f�OOO%p��c�@-,��9��Y���I�M.�2o��>�-���7�&3x�&����z�tu�Z+��r"t�A�^�+�o�Ĺ�^���y��f���Jw�Z��af��X������� �H�eN�;eە �U陔޻7�&���Д��B��AqN8`|���z��=�!�p�}�ѭ�r�y�OΞ���686�:(����P�f�. �no^�� ۥ?���ŬsV8ף�V�h� 
�Ux)����R
ڭe�}uʣs���(#�&����H2��I��@��������r��})�	dǯޚO�vӊ-O��3����e�"��q�2��B��
-�l�W'�̽��oJ���ܠ�n 2x�,b�#�8�����J�u`'�����jX�;զ�nQV�J�{��l���g�	b��Y��_��"��BOF��M���;��)BՆ�Te�H_q��#*��$���zZ���uC��� '��RZ������88%"��,L��n����;.���p��$�fl� ��
ݖ)
�Ub59��� �d�5r���n!����D��y-���
�.u���hG��	�.�� ���C-ߥ;�XU~uI۲3{����Ā�u��dsIs�Q1=i,�������1е �<6:��A�D,�s2�i������l{ppC�p���o'���O��m�Ԫ���g��^h�Z�3:�@Em���9�[m#�ܾ�!�7ٌ�ԃ�pݲQ
�S�*������p���a��p��G��ț��	)���&%��'����$W��}p��R��ji���-��|z�T����uXw��u�L�$dS�
�� OR7���{L�Ǚ�Z>v�%GS#Ť���Ә��R`S������}o�#�C{��VR?c+,w%����Uz�DB,T�3�惚��[���������-M�G!�%�����	]�t���O����q^������]d��̽�̴�N~��:��R��L#��t�b�q��%�hd$k\@��$��ց^�J�OWʕ�O�A�C0���.p��vK�ݬ�/wT)ێ�CA��b!1��$�d�g��-�?P*��b���X6�Q��P ���U;<9�\a�P�����9A����6;�o߾��]Υ�u�ɌvI]�W��9|��_�3/$�u[p�fhhh��c�l�(�| jw6�#_�������BB�O�a�N.�>� ���rb<�ں:�u�jo\���x������7v� У�����̮�e�q��`�j�c����y�'x�rw�-�~�DN��$���@ŵ�I�*��\%�^|��ߍ9�+�N����<��ہ7�y�53󁙯^:S��l�T�$/X�]6��]�H	��X��o�8��q^�H����-��rM��ngD�#�;�EE��.l�|�N�F��&�p��%�����"m7�B?�����^��j��J�.mm�������؎�5z�_.+L��^/Ư 唽�Vα�.t{�d*�o����$lҵ'��	�'j�?���x�H�y-N8pߏ3��M�XAE;Y]����(���Do���d�LG��`�7gy����Sz��*� h[%'�V;	-�3���U�$Sԍ�qͼ�o�\��59�I��U��E����$C�?p��q�ߖ���&��#ˎ�������\�3N�|�����Vƒ���	�~�����SP��h�cZs{�������E�߻�]!G����l����X�Ç����n�QQ�@|�"e��m|v,@�Л��oOݼCџM-d����|�E��S��)u�j�.$�O GEY�V��蛍�@0<��̍��iI�	E��,�k���q�E�cWdwa^�'�/�Qv�\d
���B�A�~�9ʉ�'�[��`+�='J�,�KE^���Y=sS4������{��������T�{э�������{ߓL�f������qA =�L�qe�̂�/o��	T��LK�%R�����7Wm���R�Zi�Bc��o���Og��Jze��9Q�˸�
C3�K�Us�>���K�Ѥ&;��V�����Q�JN����-�up55�&+M9�~}��a_[��BϮ��#Hk�%�~O�M�ʴX�=J߇\��-�9�հ����׊R/��'�GY~���Xj$/�Xp�m�A;� ��1+�6(�|~kssI�y}�(x4������N%8!!u�gȬ�qK����{+i���}@�>
�
�x�����\��u��A%�(�r�RO���8�;=�� ���p{�|�z\�( \	��䪕�)8��}���X[r�UL�1mxxbTH�7xy|xx8���1�t��[�V<?9>��ؗ Ȉ6g׈��? F�gce-;_m����Z?-����.t ~=~^	���=NW/��r1Z��Zu��y�~%��5@��u�`��Ä�W�gU�魹�(ⶔ[��D��E��>��ۼ{�* i?��_�f0���1 //[]�S��#�zrB¯��%���e��P<_'ŕF7[=ҖǇoK�L;�0��}�!ؤT�ss��\��[��/&��6�H�(+�b��w��GP�u#�l?i�6���D�x���j�y�m��j:ZvW�z�cQcR�rv�Z0�������Im����6���[]�]�bĜ֎2V�DZ^@}�2����E�:������iIk�z�[H��	��K�R�s3���r��|I�ly^v�ϣ�����/��Ye�Zuf���)��o=�������lai��P���o��$�/*-r�sl��7�=g[�{����@{��8S��\g�Qr�ʤ`�&�t\����#��&s��i��i�4��پ�ѹ��:�͹�d(���(a[���ElZ���@3�� ����r��8�(���󧓡��OmT���mC����^�LCכ4 �0E]N��o�	�
4A��Ȣ_�G�Y�_����I��1�G��ғ���\r��Z����7��n�Д8��E����p�u7?�I1��^���t0�ZԵ����UU��X�`}�a�������a�~,���[�>��~�-@+D�u�lB6ʯU��o���h<v��2]�V�:@���t�Ζy�܍�}�ǵ��Q��߮���,��YHI�o.��n��F���Ѿ��Ҵ���<H��j@h5�/|m��m��|���F�2�4��um*^B{&(��.��1��uɱȂW?��T�6T�,Rw�6XwzmB��	'���Go�G��D���_o_��������-LLL���ܺ��(��&�i��rj���"�yy���Y���H�~����X�{VPWwA��LJq绊�Y#@Kmn�v���l�I� n���EEG�MjA�����(\E�=��Cx$�������<�engw$�6���LF�{��vm��B�7`CS5���d�!�]�De͂�6�zS���p;t���e�v�H	�h�׳E��
����
L������N]ϕ����>�@{:�D�X�l,g�Pj�D�����ͺmPdh�"��rϊ�ě�A}�VZ��I�RKRw��R�VNb�v��۬�~8e00�Sq����)DJ�V`��W���\���j����̟M�F���!g�j;FX��k�t6S2��O �``���E�J�Uo7�Dg��}��"8u;_�.��c�,���Gø,T��;!`��t��tt�0��Ҹl��@���N����5��s=8�e[i�T�_TSSC�(Z�y�5$�Q�gN�}�7y�{51���ۃ���֒����`$���w~8�T3;d�nZD��M�?��ߠlu1��i�ΥD`�����m�����t�b���m��I 6���Y�9����Ў�htU����Q�=?^��~h�#��倮_4�)��_6�2�R�h&���@��A⮏~!���c���'I1���� ۥ�'�/�e��W�di*tLTu�YL�߭,��<̖m�:�_��ٱ��m_8K���̝�"�jFT��o����O�@��$R�����Qيe�Y��l�=Vu�Zv��C��97���)�wT������8�(�]3�)���TEq���D������C�]��9\:��|n˨�C��9�i��c����)�ҙ�È=[İ�z��ȈN=	c��a�.㣘o��:;�:��n�*���4�9�����z���8�Z�Rt*Cߑ�:�g.
�;Pq��Â�,1�.���*n������Q0x�����Om%K�H���Ir����9�3�v2IdTq�y����}?���`�.]G��z�aC����K5��n-�WLS�ٝ��)�[�Z:��l���D�*�j0��.��{���vB�X}/i�;��Wp��r�8�K��x�7��쬬�?�7�I�ۄ>~ҽ�{CO�A\كk��A-R�m��˘���v�B��R��p�ُ����9J�i�s��C��E�CDX�/W�3aea������q> 7����Q�D�v[��5mn�� ��Ov���d��H����d�y�#���_5uz��O�.sZ�Z�;�g���B�Jm1xH�rs�0
T�yN/��D�<�����n� �$�_����\O+K���:��V�.��3�G8A<gp�Y��B�eO,pk�e��5��ݤ��Zq"����MVz�[�\
۝*��О\�`I�JY#C����W#Z8�-�i�}p�ƦB/I!�������obL�f1'���O�V_~�mk�I$���;^ļ��^nL�*�A!�׍�����;)�u��z!�f|�Q��(�+�����Bġ`lRF$��ZS{<�����"���{��#��Ѭ�;�V.����@C")bc�?�37��dk��Ӡ4{++��A�/�d����q�7U��۵#�z�����?����V�~퉘���|�媀�|<�Y�is"WV9M��onn.��2*��\C��}�r�ט�~�`T�O=�M�v���d��B2MS�������=×_Y�wx���|5�t�&���<쏗xrp�K-��Pv*y�5�oTMuE*E� }#�P~O���Qc�E휄s�ݾ������B��zH���L����pGUe�"ոK�V^�q>�?��`���o7��~�Z�:�9\�11��<�W�C��D���Q����|���J�xK�M��N�ET�
��n��3DzC|ʹ��6���/��Y'���ӣ}�;��'5��A��i�3��/��
A��у(g�wѯ��>n��+YY^^���s�uֲ_�r7(Y���lQu��J$�w�7��\;���e�%��*X_��_�:)QTTĔ���^�5�z��'�/au�Ɩ���9��3٠=E�x��I�%�����V��0V����1{��� �N��T5��x�?6;J�5;l���M�w�d�aDH6�Ѱ1��|����0�γ���7���'r�'�'�r����k���U����Mԁ�6���.o`�&�����dO��P��\��	����O�����-I�����$�6@p��״8�T������ �-��p�Ϥ,QPZz������q�Pj�bK��$8���W�h�B����Z�*<ѓ6�׿eI��dD�����r��Qx�_�UD6U?f-
�`԰�@5�e���C����v�X9}@"�/�)�.�3��l3O]��Ⱦ���a-r ��7dk8��F�������(
��w$�{��C����?W@e���­�)�4%rR[��E�s�S������\U��Q��}94��ak:|l��i�2R�nC�)� ���sʗM�i�N��Krս&,bpD͕�J���Sc�A�sE��@�I"�{���&w��$���Pῠ�[���-s��v�Ɔ
�����n��hD����x���Y�v���,7�"/Q��~��i@4��D=X�Q�.�We����g{g�7�]�+g�nk�����L����XXX������ȂX��虱�;{����Wt-�z�#H9���G�Cu�6�Ni�/^��KK[U'���V|p����ek�J�v铰������Ǝ�s~����)��i�B�vո|d%�������e$�@T�jk���^����8X����ݣF">����4I_X�_P�J]�)k7vW!-B�6��� ��)Ab��O#1�/��,'�v����0N�ׂ.��e2(���n���;�#��4Y>�y�!ͱ��3��w���Q��R�'x���㠚;z��[����A�mEiX�s��V���}�nלmdj�m�]��B�vIxf|�;٦a���b�ɦ���.�}bn���0ݎ��9d���s�e&>�K�^_���C��t��NQ���b-���(�t�cH&�-j�A�i�5~���8fֶ�z�����tt���q#�� .aT!Ƽt�❨��#�aE��@E>��KKvϷM ��~&���Q��)��t8.�0�S�T� v����wX�yyy��U+k\��2vQ���=��,������g���@ ��hޞ?�
�����>�{`)��>
Lm;��b.7V��_鵹��o`GS��r�Id�pd�#���Z���r:�֝�>�+̟F)o媬1f�L���� �lM}���w_g�x���e�67��hL09և*�=T���4�x4�D�h���:c�D,F5�u#�/�܈l�J�@�Q�ʬ]#?Kf��pZ_{u�}���U�Y�c�;��3�b
�B
�'d�??"����ᡉ�QM
��=��4 ��ҙB'��n�F(8�]���!n12M��R��_�~S>���j�i�[��u�y=p��Q��S��Y��6|-<t����p�%"(�˘I���lu���z����{ok�BZF~�.B%W\�>NSPR6%�b�~.
b܇��`'�ΚcO��D-��S6:�d�Uï���gc���A:ı��<ȋ����c�q��d��vc�v�(p�Ll����^�ꈑ{���.+-Q��<搛' ��τ.x�<�p#�;�4�qNT���:R	ɉZ�"8�#,'"��QZ1_�%N)ܫ�.���J�J2�*r+x]�AX���Ӻ���׶`���s{$�~%c9�evp6�F��O8��p8]�:�Ќ'��������DS���z/:=�e���G�I����M��Kb!��^���d[��4�p�N�c�t��HR�X�aa:� �����V��v�|"u���F;�B�sK�]��lR�������Ѧ�+�.L���V����!�|y��#x*@�<x�Wj�'&p��Dp��M|�}�ÝR�ܼ��yO�d�2b�L�j�҇%�����{}0y^�D���z�z�)�2}a����E�ŀa>�)�5��]?n�<%��y��d>ƹɏ]���-<����LR#�*�Z��@R�є���Z3a���]��_�������'�|6Y� ���k��<R����P�Kv�Z��(GW��m�O����.������/m�:&����"�%C�fgg��TU�Rc�H��d�>��i4W�`���;>,PR����Y����Up�)��S��KES���t�9ݎf�c$i�rG�DO��3������ȹ�\i/�81�����k�p�U>�?�,F�,�ۦ�|y>W֯6�vk�H|�m�V��ʱg��萗���qc��9�����&x�GG7�Z��٩�8!���v=%o��Q7�b�w9ԋG����C]}.����S�Mk���.��5�l9�Z�sd)&R1��fu�y����1�C{W)��A0X>�5�c9&1�,�!�m���<��0���7�0�1g������\��!�S�����úIZ\���9�/�#u�s'Y�~�u���z�CO��`v�%�jDC�rMzm7�w���*�%;B$M��.M��:���
pQ��|)��K�Np�U�Z��x����	š�4թ�w�UK�u]4����vۿ[�ǜx�|�1@�l	қ*JJJB]ms{�c�rv�8NX���/�9����Xc���(�I��h�4�Uɇ�ќ��Q����f�-�2�R���y�"�����WMb�Y|�G$`Z� [Q��r-=�S?�������Lnř���x>bmc�mE����E�Jg`Dx�M�y²B$�&&��X������zK�_N���T����
>w է�kAI��V�v�s�6�*�!�m�f��qKbB� !�܊
SK `����6*�I)�ntI ��Q���LPWn�����;�s��m�vG���xH��.�W��|�! ��hS`�!֨��n2	��	"gԭy�p��'B���R�� ��y��Ӱ�$����X���+��v�C�qc�}�C�]x����()((�/�K�1(�tc�9u󂞉C"yǛaug��3?�/�vUECc^�?,�����rW�m��#�e(�t{l���C�	Q��')���	53���h٪�Pj�ۥlX���O�[Ɠ��uZPAM��["�=�<����E�߬U)���Q85Q�.��+��o�oDK��$�S�g������u��5���o��bwO�Ӭ���QE:�I�<�p5��B�=�6pO�R��ʒ�bSQU���#��y��ˤ�Nӡ~Nv������|�Bj��
0ʽ,�p�^7]�v6���~n�qt���lt� z��l�'��y�s���	E�t���o��i����� :�"�<�*���TU��LMMA��N;�p;dSH�Om�;C��p��nwwDD�W?`��b\]�4��N�,N5�����r6o���!��D(�P����ۃ�ou�fJ`��?�������~������+��ܿZ���L�� &Z�3�?�����6.������)�ho�2��2�*�i��#�~����.��xa��}��֗^�&��7�� ��0���=����*j���{�����l�E"�ƷC��6��ൈ�`X�'c��sx":�G�l1}����6�}ǰ�o�w��~0�nhh����{SXo��'t�OTfW��@��@�!�K�fF�Q��k��r������
Q@
m��K�V@kW���5�F��ǜ��BI����0�T��'��No:M����Һ�U�Z��A e�K�@4E
I������X �m}����ʺ�/�zo|�ο�$~�[����7��L����+�=�+Z�ՀzN�>,+d�y�Ğa|��g� .�y�3�1��T��.�ȈM<�G~���XL�Ư#=��N�hvd�rS�+~Zw�4X�F�>�P��qu����<ﮃ��~)s_��@~^��Z��p���a��MZ}��;!O==��T� ��{����:����Üf!f�B���6@H]����&��Z��wy�&8h�a�(��%�D�r����s��QFw�SӘo�,R>o�]d���T�6r�R��`	�s�"P_��>����wmf���g���]Aj5\����o���b�Oe��Ou��_wlt�,����n�qHX��+�� ר�9�����}||L����\�(�%���5Nê:�b���� ���2Ꮙ���!����| x�=��Ɣ����s<,���|���ߝ���h,���Ʀ�G/�L�}6�O�I�Tv��p�����h�#V8I���~0�&�%ۉ�<])ӈ83?���4��{��W㱱�B�P����Bf�9��swBM�]�R'�a�	F��*1�������Ѕݞ����UZ��0K@�(��q:�� a�'/@a)m>�|8�C;�����mC�q��?�Go��E)���������7e�zN��F���8��/����1Vn� ۏ��˶����o\�R�v�X8�#+�Vt�-����Ȭ(��9���'�x��Է.ti@��y�1%�_�5>�,f���8���\���c���w_�i����C(������l:p�J]���ww��͠��ڳ�e�6�m��g�b�i`�@OX���U���Xz���Ӵk��΃q��q�����n�K���\�2-�c{�x�m�'�j�w�EK7i�c�\����d� �x���عp�X�[��o�5=I35!64��$�7A4�.[�>�4�)G������z&������~w��0��WL�?3�A(q<��bE�#;�T�H���掻W��0a�B��`�^�N���_Q^���3T��0�)_�t& a�2�-������)H�o����S%!�
P��Y@��ah�Ԉ�b����bQ�>���: f�y�%#Q��(Xs���7צ��������I3���ຨ����dCޤ�9lt�*e�܌e2�i��L=��'"���u���HE��8���	|m��Ԁa��#�������=�7\V,�a��>��H0�T�=*��<͉�~��^Ѵ 3/3-���^=Q�g����N�H�M��?��X�f�c���#-����}�_%��H1�m
��O�v*T/�?��n��I,䱵��FG��
7�ų�3����Փ��ʄ����w�P�W,P���T4��.��=_FG�dR ��!�s�gNh�����;�|'��4�wxx8n���C���b*8M��l���	�"X�9&���^T��pa�!��n���r��!H?����׈���!.p$�Z�X�y����mg����Ѱ�������+�������I��M�:�ې�s�ͧDr�%�D!w�MJWG�����9��$��K^O�-�	>����_g�B�EF�U8�:2a���a9#��Y�{��
4�k1Gn�lg.Vԙ�Z��y)dA���s�����#:]�t�~����#q�����&�������c��t���eT=v{D�]�x�˓;]��;ԣO��XX�|}��Y�8T�̸�W�&st�¿��c�1�ZY��y� d�B�ߣ�1+C7��t�_��vÐ���n]�+��o��;}o���� đ��s u�L�g<�K��[;�:p�!@�T��x����T��KtEJ?cͫ겱�*���qc��4�eP��ӆܥ� �ݽ@q�A��;)�(P�)��Z��kiq+��5E��y3��|}�gw��9{�C�2���ʞ*"�p��:aC�Bg�7������{�j���}�7��X�'z�(9��B�
eK�e���7��q9C~��|MT��K��!���f|���G���T�"��v��2��W�ܜG���n@+iTq&_�23j�/㱞���3��Q��m��L���P K���;��f�К�H��%�<�#Y�ܗ�����4bмL�MG�e�����	i�VoS:�8ڨ�t⏻�����d v��yU�����RγUa�\򡎮�Ԝ�_�޷[E*_�r[;�و!tQq�.oe##%����w�#�A��� ��@N
�i�G��*#�%�f��)�,
�&)2^�'�Q��i�O�p����&9�W�cQ��a����j���J����i~(�b���'�C�s	�)�ykC}�䍢d<�OC�̚	����!iXsss8O�w���|�&
`=g��[����}p֑%Dc��{�����O����V�}}���{ܗ'�'د����<�`�h��rG@	�E�2�/�ߘ��p�g�v�.D6��ῒ�K�����s`4��Mʯ �s���-�����1YΏ�Zb5���eMl�1#W�*��~��}���:��i�/����D|?��P��+�D�R^�#��X���
����h��@�:j�Ȗ����}z�k�9zJ��?�,z�SW=���H�YL)X��8���a���M_�����&W���F�����{ǐ���/_���!w ���	x{8#���s?8O-�ζ��EA����$�a1\�A@�����;0��_�x���F���9څ���+����9�x��I6{��??�}�Y�����eşU�X��i�lY��JQ��s6���o�L;���G�o�3���xG�����5I��KĶ0!F���?M�H
�{yy�g��0�"7G�>��Ȩ�L�>a�}�~�2�6�|w�'�b��I��CL���k�2pͺ�$���N&Z�g���Hb��	���}�=Al�}���=����A-���/��z隀h.U�v������6�����[E~]e��>bљ�n'�����;����]dm�䟩5 '�+Bg:�z�,���0J:�vbc�rni2_���*�,*�i`����%)���ԟ�ة�~��{�O�-���9a��Á|s�1���	U�7���7� �P�[hM�ݥ�����;;��>|����4��q�v�:���9�y�2'��+����}QE�����;���W���Z�1�ׅ���5B^M��.�l<u�ݛ,bW=n4�J��Р*����7�������������}�	m�� .�X�h% (�6�uocm����fF*�F�]���©���=��q�U��l�N�K�y[S�Q�թ-�uDz�+�J�2�a��s+��;�X]V��a�N�q�U&2G&.o܃PZ���>�Bc)����L�}��e��4�C�9V)�*B���q�|u�=Yi����F�) �"(�@i�/җ����(��B �?L�.$6a�}u��!:;����Q8�����?�3���޸E#%�����P�q�=����R2�~�Fw��?�t
oF�ˋ!Rp�ì��⊣?���V6��Rk4�Px���qԞt`](�1ث�N?5s��9�s��:��K5T1di^KM|�s^;(��V��K�#�!E~e<H� 7J6�v��GDZ�կ,�v�V_"��	�K�j"#�����"3��X���F�9P�7�n[�E$N�}5��d ���mg�b�X�
��6���W��ek�˞*�BcҌ�)��//?��9�O�Ǿ�<�n�v,������ʆQ,./�sc�M 1�5'�+��4�3�Ш/@~}������?-�:C@k9� -�6)�u�4k�O���]��+:f#����մ�hV�����F�P�l�J�&Y�]XKcss�T�^͟��]��ƍ0r���T�11�@wa0=gܢ�6�d��S�� ɔ��]턱��P�p�%Ȕ8����ϱ�-x��9�y"Ow[�°l�kB/{�ݚ�~��i��&��C��Oy�-9i�$���j,����w �E��)@\8}Ep/�U]$7Y�m0M�%���h�Xs|����~�ą�Ԝ"H�]�1�yF��S��)��b�֎�z,�UzX�A����_@7�=6�J�����[�-�#��7���^=&_��2��ʊM�:��d�Zso�LMM�l�����O&�V�(�����Rkgy��*���  /������ՙ�[�b�9�_�;������擥'��i�}3c��%��q8�f��z���t�63��y`=�Ӓ�lq�lQ��Ts@�zz���`�D�O("�'ߜd�rRZ ��o��)��wL/�r
����|��kPu���~'��#t��m��B��e7��9�.����ާ|�.��_n+Y]�y_^{�`���Oj�o݅=ce
j�g)Rr~���m�<l�k��,R���ݖ^eo��|J��� �^E��\`ڹ��\��?1�x��^d�׿W�_+y~ͥk	�dkD_eA���80�
"�nڪ��_�嶯��Գ�ht�yK��+	H����
}"�ː�����y�`\N0����O$���:�UO����.���Km�Hz��S��AF�	�Ek]����;�����Zu����#�K�b�����f���W4��q��鴫bW�֕����|+4����Ռ#~��u/�%WZ���� ��w��"���],������$�|���2d<��cG��e�����[ڊ���h2?�-W���s`�St-R1(/ۡUa�=)�؎��kfQ��@"���k�rqU�=�r��G:o�ii����Om.}78�Li�\')v�>]��"���}|��*�<Ɯ�]�����I+�z�|�|�QmP��L///IR��$;O����|9���uێ5Lzo���F��4gj�:��]]^.�e��xX����@ J���Hl����(ٺM՜5��@j�D>�LW�K��s�q��a7����L�����L�3��qSD����nl3g���ɯ��Ee����u�q�2�a_s���l�u߀�m��������D�n`�a���xx���<��8�ǲ:�()7��� ˕l�T�[�PY���s��`��Zq�Cs��?��5A���	h�gԌ�l)U�Z���N�;�/O�䬡�!�^�+��J�Fۚ��ٟC���]μSH���A������Ј@*���%A�:�z�Ɯ�!!G"Z=S�;������"7u����������'� Y����=F�t�X�r�D�Q${���*E������� 'q݂̍~ �����\��(&j�o���@�%O9��dL&y�h��Ȥ���j8��^� ���ތ�0)�,Y��|��&x��/-'���Z�xM�
E�1Z���`_j��;чxf�Ԥ�MdfL6��M4��\#Sp8�H'�A���\\~'ߋbE�~��3�E�ջԵ��~~O_0��t�~���n��h�-(|�菧�
�.������ayo�zV�����զOw8�d0�J�h�l�"��d��yJ�}n(\?4\ϑ�h75���Т9��jz��1���:����%��R@�k\@V^i�W��N���� ��kq����N���;�mɱ�ĵ��^R�����pX�<�-� =���BѦ�6��ǋMK��qz��{� t�H��n�'�s�."G-U��B����\���>��L@�ͱ<:��!(�o���5��yV�\�_��4@�P�;æ�R�*5nJ�,V�"� o[�J�S�9v���-$*`��7V���n�oj�9�Z'��{pK2%��
/SUq��=8N���X��:�Lq
�t>}>����D%g�QY�{q$��=�rV
Ֆ��FI�Hy8^R`�1�N"���TÞ�z��pHr�2�ጨ�SHR��L)�����26 ���C2}T�C��|�^� �7�P:����Nf<?��p��������!�g��
��3@�Qh�;;�չ�����7-��M/2��G
��I��%�k@��2��rw_��̝���"��!�\3��*��"���Y��������.��>�xf�i8lX(�m1G�r�%ZV�,1>��?���V�+��*i�c ��w��+�i&�te�s�%ъl� �f,�{�L��r^蒲w��J����f�V_q����i��r ��ܣ\����|G(iMvc���W���N��Ƥu�����f�*�:�]����Z��%�����Q]i�;=m���e���Y]*��B�C��,�"�I�,�h�U��h�&mլ�iג���>�W%A��Wl�ܐuv�Po�ҹ�؎�6�<��A�0����u/A�=7Y���u���a�r���t]����8����ހ~�m�E E�{���[]�b�ʋR��+j��u�bߎ�G��I~L˟�Ġ]��Y
��6(ʐ?&n>=��l�y����/�D��+U͋lNi&_8h����j�4�:�4�Pw���<2jE?a����:�ƃ�s��p=^v�pai)�V��G(�̏*NI��3+揄D�.T���!2����Z�MP�|���{Mto�|D�Ān�7}��~̜i��p���m�;es�7��a��ZJ�#,`)��O��z ��Ō���Z}�|�T1-0��p:6}Ac)���U,�>s�>��Dz��^O��l?�C��YH��`!�^@�:�%+s{t7��ky�W��[�lvW)����||��js��v�C�lV�$n�2>��]e=���"������$��+I"	K�����
�x�'2*�46����W�Fp�
�m��Ǎ�CY�V�a�G�g��<I��XҍN��wح5RM
h"�1�$��]�o˷���߇�_:�	#�8���
ca�΢�SHo<������2���\a���2��f��[�����.�3��	ڀp5(b�pj�G9fk���O������v��,������x�p��Z����c��_����.��-f����?D��7+	���Պ��	(��Z�b��n���~ђ-Y �������9HE͢��V��A��K'$�y�ª��CƵۆ.�������p�T� T��RP&Qo��-��V��Vy��h�9y/w0�l/�j�2����|��-Н��󯗗��I�p/��0�wv��e��v1/)�?~��y�5rR9Zl:�N�V�58�,j9�_h%I `^/G�~�������p1��QH��E��zEw����+�^����K26QI���AY�X��	�'���XTs��֙Y�q~~'?{P��w�����N�.

Sա��6�۫�O�=̀:{�Q_!��g�թ���>f�/VZ{�A��F��e��x�X��n���}�[��UO|{�N��{UUNɫQ62�������t/�'p2��k��3.C�2��ۭ��v� w�e�`�.�vy�.��rj���f�yeE��<C-��޽F]~񂃒=�c�n��~g�JY�h1���o�M����<�wZ��u��u��(W jZ��[u��O���̢c!�u������v�e�9��hh���25śxE�}Aߋ?�5,\\������4B�1nT$DRV 9�Z��&\�7"	��?r������� L������ k����
0�%��i������L��/%������V䗌��a�
���A�I6��c�^|3Bx��x+$e_`g1�숧uU�\�L�|q��9�������7���q�T���~�Dt6\��\j��hq.�(ƀ�ܧ�yC��9���V��	��/^��|�K^��T�_11N��a�DiR�{���4o]�t���͌c~�Zr�r����� �S���hc�	m+}�@��9�e�k��gqU��Jp�Q��ZGd�mQ��1��ƪ����������9���Z�h�>,�)���f��B�0��'t��?ݟ����dgc�uV�R��)�O��� Q�9��l��J<^Mc�UKJh(F����h��0�2�rE����*���b��2�p�4jgS�o��,^�xR
X	���e���hy.��Gu��ſ�����nÛ�8���>�jI��k0����K ��\6��(D���@`c�qԒOg�x��W3[z�^���"�y3�|�y������|J��sqʯJ�^��c��q��'��I7�&ypk���5f=�
;����F�Զt%R�?&2����5����[p��2
��� �\���:����212윮1�|�L��[�7��e�A	�'��U0�`V���o����-�~0V�y�E}U�[�h���Mz��|�a�q�>���8G"J��#���E����S�K>����ↃHH��?
��e��y����'�&2�\���PЀ���&6��A�J�H'!=��{#q�SN��?%���=�ϝ�-kL`�<@�n.�Q2dJ��Ӭ�W@sE�	<��=om��2����;�P�T;g�����NX�7��4����%u����UtSH�nd�t�K�vyߒ��~�'l�{Þ�l��2H�/q���x�z |̓��ȵy�Ӥ�#��=����"�&�0^5ݐI~��7�{�K��G����6>��j�@�8��:�,
��l�3�ɍ*���r﯌�h��Q�_����d�"]ܸ��)G�����G������j��������Ns�Qcaވ�:dI���\t;�T����;�;�������m�Fk��z��6٧��4�{w�ꮛ���ٓ>�{:S��$�Wnd:��I둍:@'��������P���e��L7�F�gJ<�{�^էX���v
J���/G�W���_W���rC��K��r��i��o�b�rQ�ꔉ����Sܜ��B�!k�y��"|&J���c���a�&O�?�,>l�y�V�G�*�5]�>N�Ť�"c����J}�c��K	�m�j,mjj���]�1'�^�Z'���jZC@�k���
�n�c^}f	�\�W!zZIb�d�Y��l.��v3O2�/��#��F�S�G�\{P�ظЀ�"�W�oJƭ�ˇP�BB��R�����=å���8�h�!��x��}�"����;�E~�:<8[%��zB�ɧ6Fr+33W�i\&���8�$����8��;IQ��<˽ӎ�n��n����܍���>5SWW�J�¡(��_�f_B�|�z|8�IL=iOc��S����w�]�0����e�`���t{���..ٖ�R��\�Sն*���H�=�T	��6�P�5� >qT���XЍp�܇��]�G�O�>�u�]��������!��t�Y?��U��
C�]�����b(�:r��s5�8n2�x����F5��a�;~���;�[�/hk�cl��Y:i���b��h���zn�ίeK� ������)����������d�5r���6�*wbۣ_�:���6G�i�O��ͳF���}��l��2���Q�Ҙ�O!�o���q�E���7H�{��o�)���� 1Q�S�q�c�寮�*IT��8�Q ܚ��'��O���5cc�Nk���R0m���2�p�+ cB��a )���x��5liQ/�>���9��;𪑸8q���72�3�F�/$\\M�J��h����#�
c��p�Ey�+l�K�Џ�]*�EC��0�|LЊ7,6l�X�{P�q?�/�{mK��Q�L����'���~sl�LFu*��Q��}>@¬A�q���j:�r��W��7֧�6���p�d�w�Ĥ-��tS�@�͝ف�s��bN�?$�VL�@H5s�h�t��3P�&��v��'/bc��]x�i.&�|�}��Ō��+���X��Mo�qn�_[a�|0�-���dQ���*�7{�(��W|���j#1�(--E����Y���òGd��"���"�}ր�i�ۿ�n�J���vS�`��|4��P�H��P������5Ȋ���=lZ,�u����C�р;��j��5�D�}�[f��K7G�K(飅Ǒ�ˆ	��بb�R����><�+�}Z�+v'>%�%J6�g��^��|<�ﻤ��x
0�F��xn�8u��P�[j9����6M�2���I�����eA���I�$\��SsPm��1ږ�(����}�n�
Y���J[zG|	�sv�>L�s�W��X���,~�\����j��M�ó�s��%��.�q���N}Ѻ grQ�����Ȱ���,���>e�dDOȂV����}�$��Z�8�vvV��JLLL����������ҩPJJ��ܷ����x�����H�v���3�_^^��bP�q �4�A�����ȯ� ��MT�ZM���y>S�Q�B������*^HM>|h��5q3L��&�����Smua܄B!�� q�j2�EZ�Px�����*�<��aڊ�h����W@�Z�h/�N�}3�����d4'1�~��ꦪ&��w�uZM�w��y������Xѓ�604���{�����ӥ/ll�r� -XZ �y�)Ռ�9���e���}�K!H��Gc�����n�}���	Y>Tb����3�9������	�9]�W�M�@��-�V��"�WU���:�w��Q�k�i�QD����X�U���(e�j���9�W��2i�����	��������LĽ8��y������y?��J!";{qP����ү]���ܤ442��y��:p^�^�{ ����\6�M�C�E�PP$�"��!_���U^
�ஶ�ə��c��[I�� G X���uE�W*傤jז�0�c��������J�,˟qqSA�r������݊!	����2� �P�������� ����B���y�����-15��>���&�������w�Sm�>~���b#%�־��UY�aK�#*�Zn��<H�ĭ��c@ӄs^W��=p/�<f�]^�֮�u��.��{����!k%�����U���|xW��U�!�]�A����O�]Zᶅ�ײ��STT�w��.��a��<'H�f���������Y�g�L-O��m�vn�@�G�� ����S�~#�y�9��"�=]��<�����+�_�ȍ�'�	�Di���<�k��5�@?��P�d�g@�O<�a��5.&Q�{�_Yp�϶�d��}�꠯�$"��Hܾ��iO�T���@��(����,
�@�����5"Иt����J�?�(���7�ߤ$��S�5�*��7 <R��B������M�/���R�L�t����L��Î1��"Ǳ����F��6�\0?qq�EB�I�j2��u��c쁌���\M�>�F3�'B7���6������ɐ�Ֆҽ.5�'�O��}3帆f�6�1p)��g��a����=4����<���YT��uC�7{�f����&g
�WTT ��W��u�#��'s5f,���Ϻ���Hʳw�wܒ��N��Ze���%���m���싌�qV
�B($ 	(�O�痢u��L�0���%ΘJ{�����$�L����N`��K��SR	��K��v�'��,�W"����c��>5�3��
ӦG���`(EgJ��SW1T�\.<���)(8%_�L��Kg�=����p9��:M�� �f�1���M���L�����ra�O0*|��d#���m�N$�j����2����s��n6|�0*Z�-a�)Z��d,sx���0�x��OtL4f��'x�v��������0�}<s��GΦ�&.'�.��qok��+��ᵯsC},%�9�s�+��M5�"�?�4���@W�ևN�:��Lc?��3��D��|�W�x�L��J�qtq�q����Q��@%0m��@! �P����r�}|�3�[�/B&�r�NlD��K�l(E܇�@�n9}�=��Q56���@�9���1 2��t��u�E�E�E�t/z B*��>�U��D|!`��--���{�	H���!�Dz��#��p���Y�.knnF}�w+�ռ��a% ��T�v���D weE�a!1W�  [�&��Z�\!�&�����W�?p�ر���04>؟W��@OuK�GR�F����w�rS�vC2�au�]%��v�27O�:�I��w9�V�X����v�x�f`�����J�Iۚ�ۻ��4(��:m�33��}]t"�������JX����`��V�[��"*2��e�(FƷ�T�Z
����&<��&����փ%9XX��666�c�̋�+�R�+�4��' �9{)j�H
�֑��Q��I��$o�3z���q0Db��`9�����*���k|B"ѿ�^}�'�2��W[�_J�x�0R�X���A���:���	;�z-��WȉUmw���@�}�V�AZ/��I�O^�f+�]�m��������14���<E]��{��b[�!�T[��aǒM�;Ӽw�sc�Mm�t�Z�J"�1��,�C���Du>տ�c���X;CtW��2Uަ@HtpΠb����ߺ(ʫ?��x�c�/�Z1kk�㪎w2V�)D�n��� 2'�u�6���<%ل�0��]�u�՝��{�tzߝm�ES��1�w/V�Q\�E������\o�5(�4�L~/,,<u�S�p�Z�9OZq(�7�5��`��@�B�A���e~�YZ�I����?CyhC˫��#���*��J5y&�o䟋[�r��Y�m#��
ر��\���0q!m���������	����d�����"%�f�`�x<$���$��N��E��N/�+�.��V�1����b����s��A��&�q=}�p)(��@S]��G���'������8�yY)�]��Z����aa%�����#<����Ry�s���YN�2�2R�b�o�
��lM�M{z+���]򩲤����?�=���0)���A�hl(?��Y~~��c�������K��A6����@Ouk�����#s��ѹ�BY�E�!�/]�:(g�U;�%700�ƆP���%o.W3�������|p32�G��F6e%���~�|�+��1*fd>n�G����*�1�D��4�~�|���}���Lo$�e(bĪ�W���o�z\�d�!�x>�A%�",�X~pR���~R�����նJW}2�@��"�����=[��T�;)z�=?��L$��BG�$�_��G����`��ϰ�Rƙ���JE3�eF��,="�"��$(��yxaʻ����m��U�%����>���4Su~�t��U���r�����	"-&�>c��8a��sI����Y�`)\9Th����q��ާ6�z��9g\�A̶�;�tX�?�NTv����M�s����]��y��xZY�?|���&!_q;;o��vݚ~�6��nd�U@UBʐCA~0��FY�M� q�GHf�CV�D��(��o��u�ȃ���\�H"�I�5��<�CU��*ڐ/e�*K&Oj0?k6]Ơ�:^�4��+r�w�AV=t0]�H�|z�b�@�}�>&�4�6���b���;)=6U���loo�R�"�o�*��j���6�@��91l� �G���_����+H�X�|yMۚ��5�[��W��۬��H�|����&V��������)���ǽ(�]�y��Bv
��ZQLC.�p�^U�9T��(m�9�1�%�lm�A��f��A���{U��j����Uf];��+?T��~(s��sPȼΪޛW74�o�9��_����k&��}��ȯ��x8�Ih�C���A�y)�%h:��nl�rV8H�mm+�ɡa�*�oX\����Om��#�Q�,C���)@E�U�ݲ�B{����Z	W��
�c�-`��"�3WQ[	[M�-}[C����鵰0�p�3o��8)4I6�#��m��� ����ek;?�'~999������`t�\=���ݗ��r<V>���Mʅk������/ϻ�����\+�o�io}PK�<�FYV78�w�:"�����w�T�gb�������p<�1;���V��)Wk���m���ǆz�wI�԰���-�B��,��m�3)���YM�J���s��G�
m��ש������#^�8�.����L�lq��G7��QEyѬ%mmdv�����˜��o׶���d�!�W�4��a�3��:wffF�@]}".��G�@ԙ�F-]'��p���:Yo��-�}}���x�	
']ЛT�>d�d�
m�$߉�|O1���1bj��z��+�ZZ��}E��Ƨ^���J�[F��]���=9WMl}@�B��D;���,;��ݯ��o��aݣBk	�7�`G.󓭲�dV-����K����T��o|
Շ���1?�ϩ�������V;drR�e�'I2�.4w�=��t����\�6�>\�91Z7V�<J%��ց�]�������_���~��Z�:'�O��i���o�꿕J�r<�$}��Wlq��p���މj6ȍ'�6>�:���	���*�3�a�#����ۑTyaҪE]A~�����ʕ���=���n�pA���o�W�cZe�+1B��j��?�=<<|�  �c~Dɭ�Vʗ��(��2�D%k�h�bdʮg�*�75s��,��w�s��P�����<�2�s��!��;��R�&=LP��,���3�B��>z�JǇu���M�A�	z;��xA�?X�b��b�M��M��{6���z�_g��L�[�!B�ѓ^ֵ�"����馥'���������� ��R28 ��V��^GS�(�>��ݪ�r(wK�����e���i*q���k�n�<5��S�X"�V[��^���}�d�;D$�n��u빢�H�u�\�]��� p;����@���]�?���^�H���PC����J�(1��!�e��Du�>�y��NXM^��iT���;K��NZRb'Y�5����Eu�D�}��n����1�9u{<[���!¡��0�
#��k@o�Nr����1VS�tK�����4 �(@��u]|�r�f��E7^Lx� C�R�]���z�M�R�+W)�I�Q1�0H���P�`�Mkqdɦ!��`cƨ�V����ev��t�(�s�Uk�s�`���Um��6g�}�U�L���9��f;4H�ό�@��4�u}#�H����*+�̰�B���b?�MǞ��rBRp�LP?��/��7�F�Ov�zn����v@�"<��o�|��V���c������q�R]��>5\b��k3��n�z�/�R�N?l��>�.��'f�],�T����mg�ͺi�T�:s!g����&$����W���������>�k �e�?o��t�:/X�F��:CQ��l�uO�_Ɵn��.GڞWs���s�E����8��lٔ� �0������
X�'hl��Rc�cOo���~�����.II�O4�oESs1ϱ��C�#s�=5ט�`����"s@.ѐ�]#	��Iؐ�ć���u;|�0���v^nյ�����c��_9E ߸}��l��<8n!%%��r���Sˠ�����.�0���#>�9�w�m��nH)�M��11�]��%�X&&� I�lģNlnA�� w����a�uc����l��e��Z�ܻXH�h 9W�|����y�P`©z�~�B��i\�Xi(��k��ȵ�ҧ�gJ�i(�߃8έ,�w���uL{��P�����r�5���,lc$��%�,U_}�-k��ک���X����(L��U4�@.�LD�)���.y1a�l5�����[��pos�m<?�$����O�̔����&��Y���ca���t	�wY�[����άe		�[3��h�M�9:(��бA��W�5m�P��k�L��e_L�}Ԥ�S��h���_~ɴ��`���]�Y�E���_PG�����Vn�\��t�g,�#`)Or���s���x{�i1������Ξ��X��rغ�Ij��a���8jI�˵�[=�S-}������O#@�]���􋎙
�yj?�f�Y�����P�fɸz�V���v$v|��uzx%-���_���y�T1�{(�[Jx������ �k��2�//^X��Cd��C���u��Ɛ��h�p�o:1��'(�
����{����ޥ��l|������Y~������RQ$��RS�r
p�2bp�׺&�]�kƫ�660�X��עSA��� ��𖦦�<�A����!v�m����f�������ս��M�3
��B����6����� ]:�%f�2/����ʹ�Ɗr�F�t�ww#�
��N"=�l��]N�����ǧܜsB33///�Iӫ��ś>>[��IL$X�
��,�d���ywg�lf,���U1K�{�p+�Iݒ����������'Ds/�7�:��S�Y��Z Cg������KQ��e��/E�!P���ا�=ߜ���E�]g/kPƅ��q��=cC| �=��\����O���%�O��q�����R3�	����e��h����`���hx��39��ʖ��?��(D�5tw�����³���$��?u�R�{�6\�7��^�[t�2
t��;�"y��"\(����>��,ᷚ��`�Woi��!��������f�c�J��}��]�U>�G)�\�]���gj����?ɬȀ�����V#=l�}r쮧��D��>*Jp%1E��f�F'DKS�����OJ�U�o���ǂ�1ʟL� e@[s�`���2�>��NH��?�*�5�ڜ�ʩ��n.�*�����`d����6�<∘��WgܾqR^+����9�S�u�z$�nk$��_[W����!:8��2�97d�0F�� �*�	�a���b�n%��Um���x�U߅��gs�̠�5� {8{�]�l ���L�m�KS_�5{�R�N⪠D��[����}�:��t�|�!�X
b�3(2�3���ȒM��Mx570���;�/j�7x��P�S��X�zіm��!%#�R������K��M�����?���2��Q�鈫����ʇS9�z�Z}��O��(�d%[$�#ׂQf�_�3׫�G-�*�v��T�w+�
��ϐ'�#��ɸ���Y��d����%4Os����l�L�"���*!]�L(�c��xU���W��b��P�Wȕ49H�8�F��z'�{x4LL�)h%R�7h[XlȾ\��5g���Q_�G3-�ߏ������Jq�\/,,�5����Z��-A<�0���0���իm��y<�}/��\�->�24꓎.zܨ���w�Z{E��?�>��M��d�*�!G��R���nO��<L�[���dWm��q��?����/�X��	}�g.P1?d�ܩ��Vy��nؽ�B�Z3$�b����#5"��@��
�X��)�9:�.v�v@�|�=�a-}6������\ޱ��㛵�`W���|��e���b�"�s�ɯT�պ�ì�&xJي� ��o���� 
����D4l�cy���Q;d%�;�`�K����3e1H+�OS�����z,�c��G��aa��&�Z5;JvA�7���Z^7��9
�a3�+��-,P̧��R7>H-@�q�Q)�SG_���t�ˉ����q�=h����Q#�/���|�o�ɜ+E��6�}d��J
�o�Y��
�8�r��d�T�B�C3E�{Șb)�%w�e�|����)--�!z�d$ar���͎��C���V��Q�a��O�F6Zǔ �Ѥ[ٯR��o���Z���4-p��9��ꫛ�̎�|�҇��
M?|�nl��j��]�p�X�Ճ�ߪ�ɢ�0o��(���>���g������֭��P����I��i�s��&�/��������+Z�1�|`��֥���==�c�����;M�M��/F
F햝�F(	߀�~|����e����S�aKs�{جN�	i(g���^��:��|���?m��?ť 4�yc6��نƀ��_�E��[O��h����Bwq�ª�9���!������������/�bXz��Zݩk�0ju���n�2��/��b�TQ\\�!�ĳױ�Q�3�ֈ���t�%��$N8�}靠Kq�i��ׯX�S����吀2��V�����wT�	2�8׺�:��q��1M\���������R������d���gTD� b��wMa�;��B��yu-x���wM2W+���=F�i����G�&�Y>W�U=eff������5��	o���s�qlH�OD�P_�G�z�J�0p=�j�q��������E��D�9F'A[�� ���u9��ݱ?�L�0��}�au�y0&`��R�Esij��������'}j^�T���؝���n��a �O<;��M����I?�O������W;o4h?�MW�U�vgA���n����Ai�n�n����F��������z�/8��}�־c��8�S2g�����q�_(���v�ʥ�^�O�b�����e
���D2�t\��С����|��\Y_����ׯ~�/X�|���X�s��z�I�����Q&*�@~��Ku�Uc4o��Fŭ_k?>��X�k,�xn���,�pP̷��uAS�͇��V'_c��IN�*?� ��c����mm��|HsT�	���O���?N�N��m�%��;��9��ۈqZ��(�ɽ���@�:���c�>j��
UK7<�/�g�k���Aϩ����wt�C�$��s ����/La-���hw�w-����L�� O���F��8����" (��Q��C�0�1*A����-�ӂ���i����p6kdd(V6{*�TG�T�7v���j5�ek5��fRE����*�]8�����5������^�� TgD��+w��H2��#B`{�yK��������t����V w��G<���#B	�¼?�����Ƿ�s�w���lї|?��%^?���[�v�H�*�n~��yQ�Y�O�� ���	�T��A�-7�C�Q>X�%ѕэ����;s�|Ym���n-�&cdF�L�k�����%��9�k�;�ƫ�]��3ሏ&5A�(:���VDm�{��ߵɦ��:�=9ֈȉ�X���8\�P��+,� �������<���a����E+}1��m���p�,^9��������v�Os+'UO��GVQ;�B[��e����˚�m6�U�|Z�*[����TvYt�F�|I�br(U?��{����[�	���.�D�Z�u?�-��t]���=|&F���ǯq�)�`	��jh��A)_��T3�6h��x��l����0��1ͶЯ�B9m�]�^'d��p3��Ƣ"�l��zD.�Ocq��de���)�`�-����]���oL_YZPl����aj����|�SK�_�J1�ʨRlU�}��ZT�r`�r�u����6�ֈ�~�����fQ�:�z��H�%�$aEr1�/��ad��M�~�8��P�q73���Y��yK]XQ	}�)$x��'̿bF��ss��wd�T��1�A�SgzK�&0|����2�r���k'ó55R�M�����k_
�ҹ�v���^�����Y��r��M����<�S�KJJ�<�]�*�;��v��'&0�7��:��v-{����Ȫ�q5g�3v}���hD�Gp�����bU������V>5^k��!6�?1�#U�Y�{�e����=K���X����ʝ�5����s?�U�\B \�I��D=� ֑��v��љ!��~�D���%�2�.. SD��]=����Wt��@��B�e�(���YⰡ�������ͮ&���D�t�x^�����
w���UMM��i�����А�M����UF�e��5��N�x{���� ��p�\	h"��6y�J����8�C �),�+�R#1��g'���'�6[ϵ:�)V5��p7�j����m�lP�p�[|��Y���٣& 5s
h�БV��+*���?�ǟ����޷0!c���eH.�'Kڳ���V��ؑ	?�������<bڳt�.��K��t��g��y����mq9y����A)��D��Բm\q~�2��)��n�O��
�?����Zv�J2�%�L���O�ѳ�$��QD-Q�K۱����Y&'4㺄;���*%Ńu�!��u-6<��ؙ)�M� ՟m>ӻ:[(^ ����$:h�C����<���5S㠥��?Z���k.��-'�y�1Ȉ�ʶ+�~��	:�Ϩ��8N֘���'~���cI��<D0��7r�0ʌ�U �D����.��>�G�G_�#���R�n���IL������R��� %��N�]�Z��b)��P�ӟ�K�`��_�� �� �uA+�5r�9h�*?�=<"�% ��.3�1Up��6����s�eAѾ�}�k�R�
���)��W���hņG�k���\�r��_��p�M��b��QV봟P;97=�4b�\3����rR�����h׹��v�T�$m��-�\��֞��~F�V=!��$�v��S� ��@��h�<CsJD�i�d2��X|��gU(� D!E�_ѷ�M���/#��e���\�O��J
���]�'(
�$�=����A����V�_Ђ|Qh��477w44\�9-
��b<��2\��_�Y<�n��̯����o�g�W����aj�����V�&y;FU3i��.;����9��,�P� ,&�A��
ݜP=<�y��_ޯ��t5J�8y���;���h�}_�^��f�}~)��Aݩ?���p ��x�Xu��V�8��n�BkG������/wg��U�ۅ|����;��#�,i�8��H���KC�>���	g�志���5δP��v��NJ
�z��~�~�ģ�$ǐ<
��k���~���k�6�8~LN>~M����3~N�U����eՈ~��s1 �]�Ǉj}!D�8&4&�e�>����U�6	��Ji�^��eed�1���K��p<�8]cx�"�=Rd�hN��h(M���)�����'��)�5*���f��Q���,7!q����0��<$��w�8��۴��q��X	�ĸix�,��ݼ��u�}?\����v�6�ײD`%h۶�B&?퉨����	�!<
�Wy���ń�b*�iZ ��6C�����}�#�t�=Q�v��G��J}�;�����ظ����g+V�;]� C��~2j&�Hn~eb��3ײ&(Y3� ؉�K���n�.�wQ�e��|��靕��6}\ɤ��>���cH����-���QQb6Ԁ���MC�|S���:�e�
�*��{��@�"��!�B��+�5�T�!f̈́�7+��*�q ӄ�����ަ��c@����
�]@,��I6���E���������[�>���a�����O�X�^e���(7�fck�3h1�-�zs���vBLL��գ� ��c�������=�ȣ=S2:�ȅj�P����lXm���%I���$�'�;�gi�V~�rS%�.{��5ldz�Wi���2py�&Bg�nd�=y�+�z�2Z��M�	��K,R�[�����d�;Mx��}k�X��[z8�)r�ں�����o���3� ����W���Q�f�Zg6w�E����o=�y	�>��M�c�.�=���a�e�r��x��hI�^�V���W�}�.b5��(2&�Ӑz�{D��-�	�f���7���0G��,z���P�#"���⋬p"�BD�_�~=q���>�Ђs���	�V�kI��|�b�II�v��.X��Y�^�V���E�RCl�	aaIq���M��!�/&�b�'�`/�L�{G�� ���r\�T2���
���ǻyu��'�x��+q���I�2a�U| 1�V���3��l~4��U�4�:e,L�Ӗ��r'��0��ڐ��z�Q2�I�����S a�c��=a��[��K�5px���(]؉Ȣ�͵��ӛ�Pd���L��8U,x�F��i}��P6߾������v���i3�2�tyR�ΔW6�NS�����t���� 3H���㨭�ߟ�@"f�LB+�m����r���b ��n��1�߫�<�Hh���O7w�-�7���v�8����/E�$}R�Zp�L�si�s����ٱܭZ�Q#���T��Z���i|�!�L������SR�F��%��q�l����]n��ߥ�_���5$q�0ᩗ�A�nB�&Wx�����)��j��{���u��i�i����M��w�?��������|>���$���A����>�_q7?�����@�RA���4������+l��2�P�/e����&����h3n��?���������$��u"9Q״�RV}��B����cB�<�5�C��~��܅G&#�$=杫�0R9<�K�\~d�m�z(,Yt(� ���ꊢ +��_���
h���C�vm���\g��^QV���RU��?��ATHJX�W$�u}l��`Dͼy����q���K<�����S�0\��� p�z�l��STt���˕�y��m��6�
@�}㗚UB�$vn��Kv>��O�n�p���7B���H���x�Y���F �p)G�m�!J�x�hϾ�R���G|�U[��p�8-��Ǹ�F]�/B,���T=F����=M��ݩ�V����y��֮��("�����ڷ�$6BNպf����$3U�5��P�4L]�@��w���Ǫj쟌�&�!��|��p�(b]�5���71)�I�2CR~$Ѡx=��0_i��3��io��Q9���	T��K�^�}:�EW�$Ib���6����er��Iu��ѧ��<0XQ�Ts3Cm�oaP�Jz<A@�e�� 頦����Dd����$6ՠ�,g�����Z��զ�g����w
,�;�C����� ��W�0Ɂ��W�ʎA+\k<���B)z	H�/�7��U��a�����L���w=�4��F� ]E��<�Β�68P�/��i�������1$����*���X�'x����LWC�|O�
���yxiH����C2�=�un����a��K;�gLfX��IQd+ac[�cD�`�3Bf\�/�]�x����Jry.��8B�;�U�^��	E�v���.��Ê��������@�	��C�,+�"[�m�D�y�F���.���6�U�P�OzJJ�MM�Uj��Vd�s������չ�n�C:� �i�����Жtu���}oA��?��������+j
j���%��G����y����Z�� *o����[g[�hfQ�8>�v�uJ�<��|u�ć�Hz0�}�_�-�)�G.�m%[�ҳ
���#�ڥy|��hxXw�w�UH�x���l�$LM��B�N����n����#7�Kv'o�1��5�q���;�R3���}��|&�X���\�!<*)b�ȁ4ZTI-70Ŋ!�@��ѹb�^�BЎ��B�U��_�k9q7v"_-�[4	�RD� ���ϓ��Ҿ,@�sH�KZ���+daݵ~�q4��Ef^��x�嗭���b_�Ӯ當"������(��\uRI�:���h�9��KZ2�_�?!�A.�~? �5���]�>��Y��4��ma=mr~�+�ت=.%�t�+z*�#��(I(�&@	<�f�ҵ[ڹg���t_��,�s�6p^P�����VY�D�4�
�G��U�`���%�TO�Է6�%kD�s�є�O�W8Ǥ
~�F�R��&=Z?^?�^����r����
&��60��u(R}&�����M{ɺy�����K��]4��dx��k/5�}��>Z�������oR�YV�A���Ԍ��
Y�@���M��'d�����~:�km�BFK�i��h2�w{$�pyr����O)vT�W]L%��˴�����>u�z����P���P
 �N�^ �=�2&*�hCj,XH��˥E�_��B�Ӱ�
��[]dF�K��$h��E�Z��Z���,��z̒�	��t$������xAP��؟��o�iid��_��K�e8,"QK�ݏ�q;�V��m��+z���iw�n�J��'�e>�����i?���Y��_`kB{����7�k�E� ;�b��"��3d�p��/�@В�S���Ws^��fPs�\h|��\��|}�Īuzo^PP UI��Z�bv�ݑ�-��AV/��em� 7��e��J\�iIR���:�3�������#���Ez���L�B8���QO��>[\o\���.AW7E��M�l�o�?#j�_�y��5��#����Q�ʱTA�z9����M4�=����f�OJ';�ZQ�@����u��qҿ�x�c;A����l�m���yS�e�͖���`mΟ�!�߄St㩚�%H��Q�g�M����w�^M���m�a;��˱�dh:��32��b�f�[��WL��X�Fg�z":/*���#-�'�c_3��Ւ�<>I�
X���:���:��~�,��k{c�jr�>��i�V����N8��s�RO~.��.���3 �ӚmaSk���".�YF�b�m:�2*����ǀK���.2��ȶ�lr�������+�=L�S��C��=��Sy�C�w�y�Ghش ��6`n�)лaD~W~q�����Z]���k���,#Cj3��A���a&��������{8��'��V�F�k���+���Z)"�Ϝ����D�?_|%).�.���r5M�Xٯ=?&*��U���NÍ�`ɇ^`RFS�YK|����=(Y�����9_�x3����w����'�|ay��ɣ.m�e
�����<�C*�=>�,7VTT����v��!��j�2BHP<m���5��>���4�T%=�K�w��	ڿ!PVצF�������G��M�A�%2���!l��^%m;]Ҟ��/V������	�]�(��
#��d�QV<�VSb��q�����:N[6o�2#��D-!?E a�Ő]t�9F����� ���q��M[�=����Hf�ƽa����j��x�kp�OO�(V��˜�f���>J������W׺�2\����ѵ�>�gG�rv�W{7�/�R�+�EA�-Q*Aل��78���EsC��k�A�Xz��$_J1�-)��b�����$Qfl�Ҥ$�^�}�<%k5�,�0����'�"�^d|�ٍ|Y�ʭ0����A!��|�E@��H��MNϙ��ϴ�ʓ<l��3)H� �F�fN�\9�`��[�9��2կ�+����I����2��8���TWٲ_�-�|�9$�3��=���M���̵@XǸ���er�����k�ok`��őUF+����g/QOq�۸�����͊˿>W�7�� �)N¤6>�vGJ�'�nz(	?�8B%�O�Md�ƙׅ���S]�ӚT3'��Ksx�]I��m<b�2�����[����F��?!q;5pM"�!`��X:�~����+����=�wh�42�V������倧������3� Q��zA�Xϋ����������vލٹ/�����4D�S���4dg�>�9hʣ�����Ϣ���݁&�������mZ�Y8�/��#��]-���duɏ��!V��ssJ��EJI�� ̸�͛�~�F��7��]O�+s�j[<Gh����+_�*����d��k���ż`��l{��L�V�xml��>��W��
���6�/�[��wY�5O�[�iq�[�Q��]���9�i��Խ|*&*��o1>���L�i�<�sǠٌE�O�4���O2*'7g�J&�1䧂d�&Z���ʐ'�q8���|��R[���{�5ry�e-5�].��5��h}iqb<{:���U?N}�����8b���m�VXPv��eD\d�e��R�ܖ{���ҹKVe	i���~Er$⹝^�(t��R�Prŵ���Z+�k����������N��	Ge($T �'/ߞ"t�y�.x�����i�CS���]^�y��>���X�+t�m�?nc�މ��%�3X�J(��HjQ֥��k�c2��XJ� o��6��@jTP���`��O��>x��סlB8F(t�=�͉P��hh�47g=��E�A�t�	����m�-O�;T�?�2��o�Ѽ�����E��(G��x���<�'mp�W���I4���q�JU@To�Ų�SFs�\ۨn��!�ROP'4���>P+���v� U��m�A"$��+�)�	+WOW��u���P�(r�r;�{�Gt�h�B����9>��1^��I�(����(�����-��:6���$j��>b�ȱ�/�G��^�D�e���EҞk����~]�\���S\�$�N+����$x�6���#g�A�����M�j�wa&�UFC��˔P=�;��f�1�'�Qc�/j�ԍp⻵����̧���C����Ɨ/��q>����h��C��:V�T|��[>�X�2{#��}}��]��L��h�[c@���K��IͰ�Mm����!��u�<���!lzq t�q>?�c�V�@$�5����a)�xTe.��	�|�[P�og�}�Ψ�&��)�XiWV�,&]PN<(�G�)�w���VA;���K�u��R��X���h�B����_�,�pQ0��)�V�STi��<c�+�������*��h�Y�[-q�n���]�&[�̎�n���%-�1C�Iǎ�Ï�	6!���e1�
��x2�D#�y����6\#M��Y}�X���6{�W^�z1�*8p,󈺥�x[�a;���wtehnl��"�΅ߔ����ϕ�Յ��m+��E��$<�ʘ��2�`0/&���ū|�Ln�d��db.�XM���~u>��ge(�.��lWuL[�=9��xԦ&�h3���F��ڿک�3p����	ݽ�?�f�F9Og��nW8��F&�p2�o��D���NAt����	��M7G�bffn���USS���>N�J�%1 ق��`%�~53�k�"�ޞb���	�C��*��a�N3�"%�AXAw�cR#���NW��9����$�J��_�mR�{��3�VL_&��P;&Bs�O+�	���/�+���6�_�F"����Y��)s
�z<v�\�]�v~y�V��
�C�����c�T��+��Kѧ���Y%2�x��d	Q��W�j�4¨��QO�.�j�Ƚ��pa&��V�D�����&|��Vbr��4�,��1R��YVg:�$�L�ۼ%:F2��î\<D"�#̇sm���e��ug�?0LC"�T���j���ox�M>�q�1 Xy1s90tc>���4Npz�_7����دP�T�Y�*g�u"��y�%VŝV�]~�wnQ���&����,,V�.fBq�l�{�MY��ዌ�bX.�;B��[��8rH��<�~"?�R⽡ ��|_a#�e�ի�l)��&"-SKg8��|��7P^�X�܅�+ΨT�+��3[ac��W+�_�(� ���=�`7nMd=���~�}a^���q��xv�N����W�<Wyuyy�d�u�T������%q���$�a�B�_e�Z��n��f�ͱ��ʫ�ك$�"�j�{��d�ZL<+��By�]��Q�0��?�q�9�T�8\�A����:�c*F	�]��d�z��E�-F@�	 �(ہ�1�Vf��NRW�]GJ^�]Td�MK֙�)6j�]��8����O���\𯓍��*rϏZ0��N�>k�~5:^o���ڂҢ(qa��D�Nj9D�TV}���N��le��k-���/+���|«���e��{ &�ίi����r~*i�e퐨���%M��R��ω�K�����e���v��mRg�,�/��N13�IN�g�<iY__��ǧXd��2�`�|F���h 6�JǫRO¯D6�>�P��A��B��Ƭ���h��F�#C���(l�i��m�3��r��1�5Q���M}h�MAO=��g9��ʺ��a|�
P-�m���qXL��,��:�	��]�߹�lر�s�c��>�ڷ����ڇX|��w�s?J��ꆣ��4�P��//Z.�}#��\W�9�q�a�W�B����q�L����~d`f�E����+���"��AY�	�-KPHsx)E�77�aڰ|�����a���.4ߞ�O��.���� �(¦ᖝtJ-�EN��o+?^~��L'��e��w7����:��g#(�)G�s��>jUT�Aa���E�J{,��oV��O��)�J��G[�2qc���qںΉ*u��ccV��M6;�666/L7�0v_�����=/f3�Z�*D�v�^(��/�xRw
�4���v�B<�b��'lo�9�7����s�Ȥ[,mr]����T��-BGzl�ć������z�G���B�u�q��X;3�o���y�Ѐw� 
��N0�h���I|�#�`�Ů�Lb����w���8�;�b\��~�p7sa�c�D�!�P�T���<�Α�Y��@Bh�w�<R,�᥸Ѩ�B�x���]�NNN������/cv�	��m�$�v�m{Cf瓶+-N��V�	cݹ;�uu�ueB�x�P_��H{齦�N���O+3TOAP7%�E�"��Ϝqd6Ba"�~*�I*��L��q[5�?�0Cr%.��|��ߩ�:IA��/Y?��o����@p��_i�*[C�,������{���{P�ȓ͠�k*��?�?�r�Tuײ�F]�Г��>�?�#�\exn�*��<ʮ��]wr=:�^m`�84_|.�.l�ؘ��"��"������2�;���X�L�k�/>@t}.�i/�~�$�"���@�����yo�?<���hQ���r#��� T@�=ӑQ�w�gw��yKr�6�Y�n<�g��r�s�i`�/�I�/+���!3
�J"��+JEǺ�<+c�	G�'�XJ�6���b�b��w3��3a�gh�6����?�Qk�?rp~ApiŨ��.*
����T��L������ъ�/7_�|�8,�ez�dX��\L�:/����#I�����d��9s���L��A��a��ԺB8b�X�-o���]�$:*���J�~�T|@J����,i�8Ė�\�k~��7��jF|J�a���Y�D�F*f1אi�� Q#��a])CT"�m�\C,.��>��k�D�صI{����G�7�ܢ���k��٘�o/c*7n��Y�1.ٍ��).����ǟG�|�s(:� **�]g�}�:`7�^߇��v�3��ӎ+�H�
�!1������l6v�y��ѧuzP��L�Z=�M迚��:<�5eR�����z���9����G?�l�-81z�M���I��0b_����ɰ\���-�A+H�����V�u	ۯ�8]w���5��Oʳ�fkMãܑ�%�GǛ�����]�p��H�����ѯ�ɭ2������<��?x޿*Vt>�s�N�Mf�Y�8����ϟ�f�q2x�1 ?��y�<C�F�z��D�e�Uɪ ���p�į;�^߿���Z�$9�ڑ�!�� t��D8�g)1Bz�����1,�P'�f���	b�:��R�
���'W���NxE*)X��R�=f�C#TQ��/����H´��UK��O�m�i�-=5k�+�d��F���L�D�=O�E��'�z�1]ԃ�s4�O>a>Ԍ�<ܚ���X���z$W�����گ ��|��I�[�R�5F��D{�5y���	��j�nQ��aˊ�I]FЯ��C��(�?��/�| ML�|�����얥y ��g�_��g��G{��j��P�:��)�����f�)5ϼ'����A��(��G8�����;��s��H���΀�B��L���<l��we�{��^������B8b+	6��Tϗ��}�rI�����p뤮��H �<#���;����w���zO]�v�&��OcWi�~?#M=�e�����[ϣ�|9`fi�lUf��A�p����o�4��u�<�?���F}��V�o�S�~?A(Q��%���!�Y!�^ GӇ<(����j��]i&��e��m�"5���5�u N.˟�$m���G�Kc��'�BK8~zk����[�ich��-��s�`ϥ�
�,���r��Dw:?��w��KS�4�(`^�}�M���c��b���vye���"��3\�L��@L�]g��a
��H}t����y�ڝ+u�����z��K �_���uK��,P�����'�qlܽI�/2�=�%�٦�8� R�Oɨ ��@Y��m�LPt r����LRj� ��A[�x<�5:`�l�A�J�C�!s�p�G�w��Vv���g�l�����L�GJ���%zh��r���x-`�{i4 ��e�Y�������.�o����w��+\q�yO�Fe�����t������f��Np����T|�;?�N�n��BڹRж�v�q$G��Ef+#�Lf�ઽ��Kÿr#m��6a�{���s��~}fN"��?�/<,0u��>)�=[��pm����.&�ȁ���W��CÉ ��yf�{����	:�	��Ga��&��R��:����͍��5�@N�;��?~����{��;�P5����[�ֹ��R��t��N�#�&A�o���	����3WOrF��1��boh�S//��I2\��S�eם��o[�t��Q���갹��9��o&n�"+[8ȳ��H�q9Vg��rX����nr"��ɑ't]�vv�|BVصF��m���o�u�@j$.w��'��%��Y�֞DU>��d�S\��=&v&��g��x�����G��"��||�1��c��v�%�4Y	��,�+�����ʹ�⿑q��q���r�<�j�㫖���`Eލ����\nmL��˽����di�(f����2't���aB�؄���M����դ !5��簯�g7��MޤM��Y_'bM�e����ʋ�{6�&�U�5����x՜5��'fN`N�Z�x�Q@�����VU�3��_�u�G�<aiK���)�Q�:Og��MX�P]}?�;����GO�wCQ�3�Rg��dr�ޣ�82+�~��Z�Z�9a���k����i���e;�K�{��U�W�#��=eآ�}����Ɗ��HLL�R��g�C6����(cճz���p0�>���0&�@"�<�_����u6������8���qx|b�?-��6ؕC����DH��]���փ�e`�4���A���)� ����y�7"ss��[WX F�ky���$(:'U�:B�	�Ԁ8)�x*~`%�m��� +��%p�=���T����6�X<������9Ś�����p�:i���M\����ț�	y����	ޡ��&!��m(�U�p����E:R�4
]���2aX�e%�/��UW�E�2� �&3��dDt��-�;�P�%+|��.��@����n�3�,�m����KN�N3n�����p�xo���4\M8M���,��K ����q�`�����Ǫ����i��v%���Fv����JaY��ti�Q&�������ƓI�%�r�IP�������9E����џB);����\��.2|g֣F,EA{g��V\�/!7��@��π`�����k�~u�b�lG���z�#yb1L��� ��d�H�}]�h��&!s��OK�9V̉�/�=R���7cB��r@o��܉-�n��_�-���|� �
�@t#���
��x|b�I����;������*x���G����A��_D� ��������o]�+n��&����G���S���t 	����#Ȧ�V��h����_
�9ˈ�(?�接�����Ǘ5l���anǭZa�9�kl�����Ӽ|D����hS�T�nY��߳����~$�`������5~_�P����f*����z�R�����Q�8�H�Q��9:�I+=j��ښ��L�R�ѫp#�����G8X���>'�vbAv��B�߹�x���#Vse�
�N�[ݤ��{�(_��<K^�2��j�����j�FD��
2���P;���)58��QE��,��Z>w��y�;�d��B2�}{�2
�Y`��~L��f�)�SX�o]O�G�T;�]�]+�</,e�q�X��]&��&�#&�U)��ۋ�`���6-*a-��`�('/�4Y�G��߫��j`B��gY��忑��L��V�U?i&�Ɂ����  �e�9\����0�>o��yE�JJ�����5��UO=f���qq}B��s�Bp��9&c�*�8�z�+'R�c���1`:����D��ߪ�*H�'��>�;�+S��������˔��F�G�P��4�6�r˯�Ĵ
p��.�1�ɬ�XAv�ᇏ]�.�y��g�{aí��uM�11Zn�9�5�gQ��ī9>����=�C����L�&�s��'+��b�{4�8��Y�˫(
,��[�������r>;((���W�O81a���`;�=�)H��ȵTs�wT�8�d��k���틦3�q�e�η��R$�3]a� �O	|��>b�hN=P򠖍����h��q��(d@�Q���jȃ j}<GЅ�T�U�{d��櫿x�s]0������{k0V#d��T~��C	�#�z�W�s�j]�pG�\�������f����֭s�BF��N���;��E�3|������·�d�v�_׺`�]x�J��^� .��p��Rg���������O�:J�<�8�
�.Tej㦋�����*=��Q�$ϬD�u�~���MÓG�1(��Bn�n��X���aǗ*`Ɯ-��ư罽8�n��vE���� Ɵ.�<�������	&������?�������Q���x�RոO{�)�-�>�ۮ�ԇr��R"Ր�	��'��$C��H���O((&�ɰ�D�M{=ls��/n���}Q�c�1���,j�4�m�3~�N�~j[3�72Eng"T"�� R���mDO��>��R{�y\�^�RZ��*���\A�e�6ۄ�m�x��Eh(`�.hs�%L�����9 {�p�u����2�J�σp�r���2P�|Ob�|��1�s��/k��GO\����i�s�Ѧ�	�u���\o5g��Ї��n�_
]xgȳ�jzC���sx��J�=�/�T�L�w��rx�ٞ6G�~)xTN�Pש�Q��L��Z�Y��hS��$�+3Oe�*엿&�d���e1����Skn^!k��tƄcK���qd��Df�Q]o�@SAV-��0��]�*ou��a�w��/rl��==~�<KJ�ʄ�9��b��m�QW�~TL�
,��7��j����''��"��\݃J.��Q
^FX�ѐ�����%��e���}���ak?-�w��"N� �g��z>��,��_-���� P7L���k�r�oh���>�/�)t�*E�u�C��+��Vd#��q�n7;7w���<E����ch\�F��Ԝ˪��Œ>�W�WM�6��wމ~`�����P���F�=�^�!���?�U��z�a�y�Y�dqD��A[3M&��.�⳵r�gûD"�4�38�#;O��l&�l	�&��H��;fHS(ه�/q��C����J�S�U6��3��E�9�}U�Y�b99J�ѰqN���O���Z���TV�N��&�w��-������m�3!/��p}	����+���	�����_M{�(e��x�kl��L��_�6��%�A���'�mtz�����C�rz�W�H:F�[�l*^Dnn�Q�t�I���%>�)���L����q����"M;��rGZ�ĩ���>7+v�s�lj%K�IN�'e��H�3��B�Ϗw.�<<.��Z8�8�(��R��}��Ȃ��B�\(�9����a��w�XYGT��^Ɉy���Ŝ�ϓ��6��#�L{j��������|9����	J�RS<!���F����}?\�����SY�u��;qi/˴��<zk*�?S�M�z�eϒ�f�> �,'��;pF�M%��&-�����xh��i���G$�ܾ��Ja��|G��(x;�1���j=a�v�}N����а�M�H�'��z�3�y�U���<����[�&�������2aIF���8Ibf�¯���O$\Q��Oc��w'd�L:��Z]�p�u���j��Q��M#~Wb\y>B�Xi���̌�St�s����"p�{�Q�����xA�Zj�"p l��=(�P�0��M�,��꿹��7[ƅ����')dp׈���	2x�u m0y��}�Nv�����V�%��h�����hr�s��
Ʈ T�����b��m;Q�ϗ/h��7xP}+O��Wt��b���A,�|{�?8ꭁY�s�-jG4�~�d[s��WU�N�ٶ��QE񚴦n��{��'�Ob�妉�>$AF���	��_N�k��IJ������j� �pp�`2�KwK��Z�~���i��D)�� [K�J�g�*|������n=����Ғ�r�"�M�O�ˣ�j]�@6K̎' ݱ\&�|�q��T��������SEO��bV���-E�A��85g-������6��}�����]��;}ts�s\�=���em�ք_k EOM�ٯ^�I���ٙ;�R�<��#�hQ�7�۩+u[�g)�/e�F�9�Yă��J�����X��鼜�'y�T��ߎw{q�5A����O(����hb3=��/j�=�F�F:�$�k87�S�����Y�G����j��h)R܊�wwy�ww�8(-n��ݭ�Cq��{����;�=3��L�쳗Lv��k5Y������,*���KD�׊7'WH�v:���u�ci��dY���I	$_V&��/Ĭ8Ss���3@�@��8�*E�V�͂,*�_���AT�+���~��;��E���$�~{kb;,����m�;�s>*.�����k���8S���F͐�T̄ß���@�ݰ�a�1PKEV���0SO\��B�O(�9)��>^�H(�X��P"�%��B$�-Ի��B���k<�!5�s/!�Ǧ�g��v��h$��i��L�GN�;h����j_ydt�ZZQZI:��S��C^�=���5��)c�
F\���2_>�̋�V,.�Q�1G��[�<\��_�Q�'R6�+}d��_�Y���B댻/��u��S���s�� �p�rF�~�9nͅ/�v���&��na�Ԗ���D$��h�O�Je����>�o[��zm:�l����h7	"��"J9:�Tw����|�X�1�+V�͒K�1$������"�~�}X�ryy��A�_9��ﴬ��N��?��x��$ f	~�>n�'�&�aT�#�x'���:�y�$����kri�{��6_ͩ;{�x�9^�,�sK�ھ^g�b:o3�!7\�}Mf:��|�׫�w�r���	�t���!���y���	:��K�G���S n��oY/���V�Tm�_^�E�h��D��1Bؼ#* U>�i�R3���Ij	�l��qϲ��>vMw5�喇�q1:"�c&7_���1���f\'%BY������u��^�͞�w� ��Ƕ�֦=K��g��+��jpk#
�
��~��	]�)�N�K�����' �q)�du�0X�� =�*�������
���R��B�)։��	FJGU�L{����(�a����Û�H�	�Eм��vO�T���1��>	�oy\��u�F��
�?���mD�wO=�{�U�����`�:oy�`�XD�{��+<�󼳯^�Ԏ$-w�^���ާ� �Z���w'�ߜG������_~`�t�H��{Z�}f�K�<C�E𖹺��#)�6�m��M���!��b�+SC�`���N����7v������w�[?�D�����2Z,����w�/�S%��f���S��M�#�p~��2�U��F�.#���|�Af�����}�߱T����L�kW����wQ�3U^M$�`���XG�#o�V��~q�AǩR����=a*���鋆aq��u}=55�~�5,X��#z�L�I���ǗJ���IgSS�0�ϻyf�^�� T�χ	6����`bKUCFD�Uu���z�#�&����맢[H�T����P&y�л!*?���Z�K[�д�,_���w���P��'�Z��NĴ\V u��'�(��n[���:�Q��˖�51����|��W�Dw�����2����:��ŕ��%!p�қ*q]⼺m;ӡ��Ӵ��H.$&�q�RE*캫���r�He��-��%��/D,\�+��~�H����K�@���
y1����DGtϩ���=�� ��.8.�^��];��H'CQQqX����^�1��ߙϫZؠn�UP��Q��?�iM6�ׁ�3U��HW���x�t��wL���1�6f�nģ����rSKѴ��5"�9d]O_a*?ژ1�ܷ��.4��.!#|d�X>���c^��ag �G�?�� �'�t�'�3Ӭ�gB�b��.�R5W�ݵ�3�����1L�p�~ǖ�$Geчݥ7(��5J��2�k�}/�F��:"���Næ�p5ǀ/9����߫���!
M��M[V;ͳ�ct��
��6��Læ����B���߅��Z�0v�R㳴4Tlffn�!AV�X˥�}����ǉ	`k��Wpj��'|r�M���CT¡ꢰ�_k�ᕡ�f�ǜ�iZ�!�CC�q�;���9_?!j�U��0�C��#~0zyZ��p��9^�bZ:.$��]\<`]��9��j��+���!UE�JE�Ό��@1��9����#�/�y��pv`wc���C�tg�쁷-E�H�a�認%��7!r�@)�}���q4Mi�����2��8��p�o�ۄ	;�.L���?�D��6X�	j��df�B�	�)К�A�4�F�z��1�x7�~x��O�Nh��.��N��9���ƶ��ʫ;m�e�)�"��?��$�m�%0K��7g��[ ��T.x¿�Su�B)]�~9�B	��R���h�m��������<r���)���<$����K�c���A��R? r�m�ˏ�*��%s�
������|GC�9fF���h�}�^7�f��1�.������y�����[����V�e��<��(l���<.��ҝ�.\������p�ꉃX��`��!:V�rk;#����Sa'�zin�2��n�p���]?�1�����zZ:.4"<"�R�w�=��>�)l�����ya�Y�/T�j���A{v$��I�����ѲME���Lbߨ!z��Dߨ�F�[����
���sB��u_��b����|g��֮N/�����I,B\��ӕ��E�7#͔#��
'��jK1h���O�{˦��z�ǡ���p� }�2���2
��M���,)>�>b^<~�]�ݚ�l���Y{<z
^И�
~S�k�Ʃ�ta�c9y�����W!��fʱ�b���<�ƿ5���O�����9�;�Q3K���s�L�!�a�":��3[�JZ�;7��H)��m%|�	 qD��-�S�~�ωJ!�P t�(���;lOJ�?�1�%*��2|�q�;���l����+�5k^0���ȷ,���O�-�z���W������Xm�nYE̾rJdw�V����~1�e�y�c�S��;�S\<g��?����
�c��z�r����@�ƒ����D�1pr�߰�1Y��*���_�N}s|��z�W������>�Q]Ƭ�Z�����LoJYx���g���.��٬�L�ӸSl*ŀ4`�W�/>�w���2m�ӿ�Z�~~w�g�y�\քc�b��o������+�y���r>"?�L��DO{�T��*�+��w��.�2�o�ڐ?�c���&�!.n�J����=��"�����K�0���7L�����FQ́��4[gD���?�r@&����~�L��~�w"C��4�8p�L�j��tSn�Y�v8]L?�^���f0BO�U�����z���G�Yն/��� s��q;\�3�kq��w*�ǯ�����4$��9Ry���jݪ�-�o�Nm�e�gt��:��|:Pd6�u	C�2d2�F_�p�����',q���t��'T�R��MJT4z1Ӭ�;m����RˊY���k'��x9�?8�����댒y�����	�n|�\��~J�r�������L�lԱ�(!v�X��!��(��Qo>��{����%���z�����.K��,�����͋�3���j<����K2�#�r�R����H,3�޳e$� m�A�ʫ�>,u��
b=��y�"Y�Fyyx�n�	b(r69�1}=޻�����r)��~M��k�^N8@�yN�=���VV t�.�ݜW�&T�1k�����t��& &�H𫫤w_3� Q4�4�%%%�ק;���,���k���Ǯ��3���N����;hՇ�Ck�@)�Y�#i�7]��e>3[${��KV����u��q'q��,}>�I�ז�"u�$"�a�N[so7���Ҹ��\5}
�.������VL�ɸ����5]�=O3L���UV6��h��,��	�������$�F;�c��˴Scq����A����-U9����k&���L�PN˾�N��h����#��R��@|"�����v�\r�^���x
�Ζ���\��n�@��A�_GP�!D9m6y?UO �=�\���0Lh��B��,Co5�D�)b������g�W�i��r�蔻�/�3�0��p&�o�t�/�����K�E~Q�1Lb�!a$V������,}����$l����H@@G�Lb��J"��Z.��ynb�����lW�k,��<��X�Y3*��Y�=g�3��n�rC��� w������c��7�ʥ��켕���0����Գ
���L�Iڣ�Ou�j�]���'�6��~k��#�B��Ov-F�Ir��s�9HH��}�5�rٖl��)p>��iWs�Ɔ��xu[;~͂*A��,�8[�3]#���Y�H[��������U Kh
)I3r��D����evv�[S{�m�d�^�u�TlM�!�@���A��/�φEڲ��G��A��h��H�"���ދf�M�����7�du6ܳ�����0���S���O��*�knR˩n����j�����~%S�A?&�m%$Wnv��7w��s��N�ZK����X�:݉�yܝIT'%!����_�9tmQoS��6+����x1���7�wm�}��V`!����E<P�r�����?���)�;�2�~��p�����)꡿(�WT�6g��b����Q�bmjǸ�c�C��$m{:u��kw3� �o�,�u�!�o�Bbn�n����~�kc����� �1����^G��7urk���_/����W����
�	�V7^��{y��P��E����&B�/l�}���o�g�Fܛ�$L⿅�~�w������\�'���ha���<ڗ�]������nڼ\4�H�F�F����{���-ӱp�$������%w� �+�/q��"��1��Ǵ��o�l埝
8o.�� �!'���nt��38����<��߻�Ú|�VR�����o�s�g	���`�=���./�������}����9�
�n�u.DT��P|#�Es׿��u��SN�/n�>\��=�Ykjk����'�ϱ�T���Q�}�cDw���Y�{L���\�����/Z� f���`��'
�v�é�M�wտa>��ۆ�w"������I�Tnw�aG4�H�$+���F���N~N��S�l��x� &D���H�ll���L:5�s�k��4�n"н�@�n9����e� ���_������O%��2�Pqċ����� ���ܟ'����7QQI~9�Ы45	���,��q.��=��"��.��`dL$F;�pQ�� t8,4 �zT���$�ȷ0��A¬�;Ӓ-b�*��&v��	�â|٬�:���:v���=�������ڷVj���ưg�?7> !�+��Z84!>�s�8�ɐ��B��s�7��N���dߨ���f�+���d��KVf��o֖��#,}F�~��q�l=k�!D>?��ϗ�Fsv?�N�Isg*��}�.(��cd��e,��j���'Q�;�#��#=-�Y�W�'r�n��Է���,�~�O3��˜e������=���ub'رBb�o32&<�����K�hj�P�ZLz�#,�}��=�o����G)P�B���a�g�Dr)�r�_��mF�G���S���r(����Ȩ��Ң�,�U��������[���`%��giudv��cq��b���"�5�u��ys�p��y�+�*>���y�f�-�ǚP٫(R٤����Tv�/���p��5�.�TCE?���ƫ	8rܟžc4�槠�Rk_4�K�*��w�d#�3����?|G[p�!J�	�>Ҍ��04�Z�'�J��V]��׍E,8T��>�Q�<=��;�&s_�#_�|���\�����`��V�]�l�*���^�F�{�.�Lp���˦�n$L�i��%���pܹ��"ܘYu⠝�a�r�~�������'//���|�	�����.�3o3������I��j���V��V͌��c�qzWm���6g���&S�n�Ĉ1��#�:�O$��܀��]�z�6)��An��'��x��w�oo$
z��i��d4�޼�q���ʤ��h�#�b�.���7�>�ϸ�E�\b�/����\ks}�؊���G��)�.����O3��X���Z��w��F��={�#��d�i�vl ��P�h7�W44�R�%G:�5�p]�;��Zy�����HB��MZ�	��6\�P��b0�[G���_>)�Kl�#�<��բ��2����U�<N�ڶ�j�a�a���/Q`OW�y�Q�5G�g����0Q
w33�b�'��X{aޑ��ٻ�. �M)�2�����A>�%'�'-Qͷ����[�����4���0�(T��c<x���e#T���6�OWh����������\u]��r2��5:���B�F�9��	�V��E�F��i@yy��B��$��)E����oE����I�2���ڄ������&S$$'�E��7+�j�H+�*�)A�\���g��0٨.�K/N���Q���UBWb�f��}/��N���~V/?@&����"�(}�{�c�Yh�7�G1k�)�R�鰾�� �(���vp�P94���FZ�A���m�����f��j[9�S�D
N`�+�)���Aн�{/1�X���VAѡCW��t��o�n�����a���L�m��r#C��w����q�@���z@/���LXA�Ji�b�TԠ��	;�sa�@H��p��!ܚ��|f�l�!�xa�����o4�nd-z���!^VP�����"?.�b��Ho���j�|뚲��I�N�}��2�y�0�c��H�hc�/MU%5*ǌ=�^����7K#���#r��!2d+[PސOyh ���0u�	�����j#H��KK���IvȺ���e���9�o��Y�>K�v���[g1LKK���l+�9��q�@����*/��^}F#��+VKF�{&�a��I�7<{����Ч�����	�[|y���?(��h��Zj�A��_�H���.?j�����U������k/Q�T�{3�GF4�ƣ�6�q��4c��i�N�gܺ����\��T�����d=��7�U�f�:�	e0ˍ��|-bGgS�l��0��Y�k�l�S0�Gƺa/`Ƕ����S�ܒ�J)`��֣��^|N��&p�q�x��(]Q�U�����b
��la439q������he�P뗤����H�aO+���ҋn*i�s���Uv�`j��9E��,$0!�=��{ad��V�����;�&sMx�Q���t�/�	����M�A�����/��\�»v����C�n���Bw�w�=�D�$1�X����^�\iH�s��3l�4R��P�L� ��4����4��6L%ʗ����F_C��g����&{�=���c�	��X[v��ƚ|6������~��]��`t7a&�b>�QExX�E�����<F�ў���P�@0�{L�$pD'�����}�ݶ�/�C���7/=I�)��[�2��?W����=��	�/]���y}�&��3U�?4��d$5�w�鉙Å.�t�Z��"K;Z�G���3F�9~	cWM�Y�^���{���3�I�:��	]$^ց�F	;ݐ�02��6Y)�פ��}�W+���������h��;�~�=¿��6i�F(�Gg�jV�E�F9�9Bs��گ�&��ʷ<Kxn��I�:xhW�m���]�����$�=��S7a�ݷVr6���w��	�[:�����5�7�'gM�)D�1B=��I����.�٬jH�v��<��3�"�����e������*�7�6��|�[=�dL\n�ɱ�*�/�ƀ� ����D��Ť�ԅ�[-����M �j��D�f X��ۗ1=�8�,�s�L�����?G�l`��{����d&sBVO�����^�E�X*"���b/	fvK�C��Ki����G����A$�K,� u�:G��<՘�F	���� "�Bv��fq�H���G��7��]kLD�n"|�����q�]&��P��ݔ�m�e�\�
j����үg�T�Ԥ�(�qa�u�ޛKz9�P��&���[�!�\ك�������/+�o��h���xm�����JT�2\��;}!,گ�j������^�x5��ϡ��H0+�?b�>������I`>���[��ʗ���/A�O=.��2M�^�U�
Ń#�)��u-\6d�8���Z@���f e0!�T;�XLT�B �O�k���B9gCK���'m;�BY��}/im����K�{�(p�G�f�P��v��A��DTLTJ����w��:Ϭ{S��Q SIj�H/OwM�Ԅp�]�{�����Ȁ�1��QO���aױ}p�r�W�w?�"�?)��~>���k�i^`��`�����n~e��C��e5�Ȼ�l��#�}?i� 5�$�����b���X4�"��,'~�Hb�a���e��e5�/�>�x�ݟ�ZV����Fuy���k�����'��~�~jC�����ZF��~��@C����n��%�\;�m��Z�U�,5�jn^���<i�����ou�3�j��7:�RamX���{�%M���]�:��l����i,�
sI���s����m.B�`Wl�	��ך�gX�n�k�E�����)Γ=Isx�����,�D������c��u���q?Yu�ց��Xǁ>�J��r#�g�2��ee��-�����#�Jg&�hW��d��J�Yl���F�3)�œ�җ�wƬm���	K����I�_���� MOV���,���E�૲0�6X��'at-�<#|=h��NS���R��u2v��̖g\�c�|�g������c�]+^g%->���e��O������Dˠ����¤��}eI�����%w�ny�7���e��<Cؤ�]./��[$Rm�ߨ|�G����p�^:K��d��C��(�L�u�! �z�O���d���p��Uhr�	���ќ�0-$�2�%׋��C��X�NG�Q&b�#�|����I��'+)W���ɇI�S�}�:��Ѫ��pMD��|�Nǡ�I�<�ox�Ww��Wj��Q�}�8VJ�R�i��8�b����|���^���^�py[1��s�b�����	������X�%�I��;�U;%j�n�?�a�QKG���3���9��,GG�@�~Cߙ�(���=کUyɻU�nC�싗�Õ�3L��o������IQ���i{~xM�h�O�F���-%Q��X�Aм�!���{M2=X���G�3L`��;`1cR9���NǔtƐ��d�*|�c�p�=�Z�_(>!�|P���ˑvW�yD��K�^e�z��[!��:�+;;a�����?�8}S�F�-�j?�;���F��.�S$T��93/+�`ġ.S���<��^3H�;���� �r?7���5l֋��u�1zɟHH�q��k!2�ܺ4�%u>u=���A�ˌ��]�|�'�9�}�[�01X�"�3���A�r�z���5�q�����UV4�"ƣ`:G_F㏘�v��c���cL�c��c.�t���뾦�I�D�r[h��~q�a�;TQB=���Ĝ��x�/c�<v'$�
���[_�Ƹ&��B����V�yB����!�>hF3 ���m*�L׀Ӧv�'C���߸�psV<*z~����yw,��ֱA�R��}�8?Z�H��4��Z,�Pf��Ҝ$�<�o�p��.xY��V�!�O��� )n��{4D=�6�_?�Lk9�!�r��g@�ݤ�A�9�c/̏)W��l��N�XMٔ�S-qU[�_f�$�E����K��k.\Og����N'�����S2�~|�Ñ����l�Ͽ5~գ��2 2}b�Kġo��|VK����Y�&���C��h���u��+�$E��S��6��N��j����V/�?���V6��/p����.}#��N��mn��l%���jjqt�-�ʌ1k�����S�-~�Z� K���ŉ�7ݑ�V�*��$������֯prعLѠ#��{���_����N��EQ�yiegR�2�;��Y�w�?C09ș�P�F�
91�<��[P�`�6�C���q4N{m�$�~�,#�w�:����u�Ɲ��js��;�5wXnk�Vl���gAt�O����*�����0}V�"��i&��<��*5�����]�<��~L=���>X�;^��R�=�Q�?�뇙y�m�sB���<70~}\�1�c3%��X�i��U E_2�L��d�1�����D�	q�%}��M�fϙ�w�GZ�5���^2��}#����
�Р��6Eg��=^Y��I���f��׼�zZ�G��zƺʰ�Y��������jy�������̆��ڑlh��@�����V1��^�%��qL�6m��;y/3)�km�>�w]e��Ɛ%��!B��-E�m|�iqqq+���l�K�/�A�0]��v�+��������ݏJfw�o-�N�.V��}��[֮J�( 氎Y��������c&W���xr��l����/����ɪ��e��ˉ��g��d�U�l�H�F\����CFи��:��ޝ4����+p:�W[Ol��&$J��<:4$�P�G��V.��\M����	�ff!f2
-�t�rU��R�E�m��
�c��\��ߢ$5<�4��HV>初�:e�a�d6U��0ʾ�A��C�5q�]m r���ؓONs�Ѵ��*�_�O{��8�0;�t��7�0������)h	N��t�0&ku$E��IV�	��;�]D��;��i	7�����,�������a� �N�����Κ7*@�	�>�⡝�4�x1:�H��:�~3�_����s������x�y�7ªS���wyy�z�Q�#�ka\���{��?.�V`��b��¬ߦ����5V�̩��!M��{gu�HY��y[e���/���DQ~����|Vf{C���xO��|1h�5w�Tc�6JhD$����&0:�d�VS�͏�:5�v�^٧Afۗ�Cԓ
Bnl��^�W1а�]f|w�K낕-��G00�4@�1�"��%V���&����g:\�w����sl�,�{�"Dj�!A���Q����s����۫�5[��p�!�lzԅ~���P}��PHer5�J�sLE3&1���\,��_���m4��gn�{-�tL,;��*��r���\^ǰ��ݹI���g���K� *ެ�x��H����d;7�uã������w)����9�7���� �[���a��#������Ԟ�Y>C�';a%�qJ����k?�=\8���m#���dd��l�����]�,+��Pl_�� _煫���93!zBRRQ&y�=�v��[oF�����^��<#&���: ��8���9h�oH���ߋ}��N*)�@��ۅB<+��,������[�x���(���u~#��a�R�j
��X���]c-0F���Pe��keZ�ϱ��Ձ�y
�����[�w�� �#�'a�8O�7ϋ��}�ⷫ��lLHN����i���fk�4�ӿ8�J?�YKȥT;>
�ܫ�QQz���&��%��0y����H<�[]�͑����H+Oy%�7���o3���jv¤�A']�h��B��.d�� x�� Z65�ݶ��5Ɋ;֬K��i����5�N�Q9�搈ƿj�!�+}��n�����׽��Ie�w���N_��;���2�}w�ڜ��?,�)^q;q�]�?6��X��.�K��l"��e���s@�u�#�2I�%�{�%����P'�VĐ���ӵ66�o����mL�\��I�����7�N��7٪�yh/)�'�L鋽�+�c�u������r���̕�X{kF�l��?��Z-h��V�=�Ȑ��y�l�b���Ӑ!��2j�Ĳ"�|	 ��Z�6�l[���t��0���"�;�2U|���w.2�W9X���9)��[�"@��ߋ�!�B�?P(J��N۔7ި�#�)���[���a� D��������}�9��w{T�A)�ݳ��� &�e����,0�c�!>���8<A;"��"�8H�O�h"�8vҲ@��Ԓ.�_�I� ���B�M�K��5�J�]�	����gmG9`�e1�&�Z����̅J�==�(hvo��'ϩz�:hca���C#.ݴ�*{�є��>S+�Rn<��F��ۛ!?X�������DAӨ�td.����G�kr�|���7��vX�٢ý�SW�%F��a���m����fN��%�]-]���"`;���Z÷"�>��k��4,�ǈ ���}�����{{{�@�f̄wb�l��];.D<c�f���~��V��	s��
~���:��O[C��g/�lJ~�x�Σ/ivU��+���l]T�������&�"[�������3l�p�vU��s�U	��[�h�7��.�`��*1v��I��ti|�����m�N����T?���^����:�.�k��Ť'��n�IX�B����%��	�ݴv"&#��JL�A!㣡��LL�O��\��w��[|!�nd�hWxɷ`�h[��h�ޠ�c�9�nm�M]#���jؒ�9���,�������'��_��%B��ݛ��g���Z�Q��|܋�\��`N5銠,wd����F�)caq���A�m�߁T}r̃<�s�An}����1�u ��w�S3�=�ީY�K]����E�K,�N&�D��?�O�Y�b�,|G�f�e5�6߭���)������e���x)$��m�����f1\Eӝ��;��[%�8�[��>�j�ڋ�&|��f��v0i�d�ty222�:�+<kP��(��s���� � �fL��XqÇg��PT_�I�u�����G�Dv�������Q�������Q8G�
8-���G\-;�yM���?��A������~�����h���.3_�l!!g����H��/�gi>�}���*R+��` �`�&li�	�I�~	����X�AQ�1A���խpEí��W���|5�֥>��W�n���p�x�={x74��͇A��"_Rl�455u��`2w�~B�I��[md���մ<�V�ׅ7��98�&�>CԿܱ��ք�f�L�.�ѐ��[֧[��y����%����f���L�WTT�I�n�O�i��GtT�b=��F��q��\I���W�m�"�qm���v�O��� �/��� ��) ��E��n�4�� ���������p8��}��A��l��r%�-����� (Y%��x��Z�
��Ƥ�E����0D�*��lT9�ꊅ=W�%BA��;�M�xԂ��O���'�>%�J��~V3G`iH@�v�i,��t#Y�'���"	}��_���,�a���7�jF���'.��Vy�P����_O�G��t�$<�z���R�*C,��պ
�$�^M&���4��n�����йb]mƟ����j�k9\��)�z+po <��C=Ľ`���+,*�W���$,�&�$hb����@��F	W���Z�6��@Of���W�G�0r�5�d\��s�9����Iݏp�T�3l'�44���]<��B�wg�:�ߒ����D�J�|��-�А���ʫ�+��.v�vi�Hu�j����Vk�q��R�W�q���Y�謹�F�:pø�������s�r4�������]&��jLp+䜧��F�lQ��tK��5��Ș�PL���w���I!�K����7�n,�7����+���T�w=Ę��"H�ڑݒMi�S�x���m?��q��,�6�nŸy�BB�oNK�,��E�[%��@f��I��ޅ@�V�Rr\�����3.1��J�*��d�~�L�H�0l:��/�_&P�c��H�K��~?�Y��ђ���`��g��"�8阡�s��t��s{�o��t�ħ��U�C<G ��<�_����sd�$#��@����Ћ ���u&fZj���>*�b~sQuz�7���=BO@�[!(������8��#��4��K��hW+&'P{k�Z	%
=J:7���'�J�����_�7\&lI�`�nq���`� ����-ӄ��GŰ1�R|����Y �Z� �\d|�~�>F ^N��L�V����z�7�฽�S�=ֻ���W��"���>w�O;߹�wg�@�nݐ6n��;c��(�9�q��J��<��k\)x)X�X���y��||Y���9�@����Z��ܶ�G���֯�"�Y��#zQ+.�
�����tjd��f�vo/��af<mD#��d��tW!޴�e*�yx��X�j�6�"&���\��1B2T
R�"�mAZg��UL��e��b�Y�����t�N뉬��݇��n,�2-LK�w��T7�>���a��d�rB�<	�jv���n�����F����὿�.�\�ݥ���6��������k2�~c�ّDFM-<�4�vP@��Orv��C���?&�r����J�������(wС��!p�Kn+	!�L��>����.��'y�AQ6
�f�ݚ������������@X�_P�sXP�M��|�/N��%u`���kj��q�cߧ�K :+F�y/:�ڨ��(fp���m��R���Y�g�;�����c�Q��Ğkg�V�#�ou�|��'�[���+�/�i3��x��(����+p�ȴH�n�Sl�f3Y��<;d�9�/�E�m<Li��$C�.��^=.jf���"`̛�ie�P|5:�����!���n��yP,ա��~#��m����/���A�8��Y���z�	���������s;QV%"���1^��W��]V�bv�h���������E8���"L�G��|k�"�	31�9?K��ɷ�^ʐ�y�|ͪ�u�\
�qh�+TKf���#S�㿃��lOX��m/�9|��c1Wm���w"4qʩ��Ӏ	�;�7�D@�O_.�|�������ov��0	�Z��^z9����]ʍ�w��I�Pt�2'�-֘����t����D	�sx�u�Y�6��8-/��F$����*>��5���%���?c�U�Nգ��q�H|��r�z� �gQ�wC�D^w�1�d<���H:u��N��P����+��(\�ZOP����u�f��F���%���f;�A��,}�V4���pɥ�����-�����yq��ޗ3(�#m>�DC�[��>9�}z��j�d�*�}'`����	�h�T�G��E���"��ַ�9w� �𶕫i�E�,�LO����\o[d��F/�g��"=`���\H7hY�2z��@+,R�`׿�O~���B�J�.Ѐ��d�?�7 �}<��6E*��*��ľ���}��U��tV t�«���x���fk0Dҥ:�:rF��<�轗��XQ�^{L��l犵�����9`��*�Z�֍3��ٰ�Hn�}�s}��5{��^��ߣ;w�.PX���6�c��9}��u�]�3�zCD���J�3%�*s��x��R?N

��q��ȕ��hA"��=O �<��N�N��i� A*w.]��l�1e��zON�/	ʀV⢔�ۘJ��#!��XL̶L�F��~�S�b���R^�˧p]}��^�c�LL����

���֦�+�0�HZ��V.u_A&�/��N�k^���oZh3q��P�ކ֓��!������k�H�sXv\�F�}��%Z��Ǜ�q���	�~tu�'���?�XC���7���!���qO��D�^L��1\vbc#�K��HC�uH����D�wfdq�*��w�*���:��b�h���y���k�9���=����`�Q��?X__��>I3�6������镏���0�+>׳ݱ���*�ɦ8���ʨ���(Y�@-����:r�-�س;��y���=�LS�H�������\ٞ��62��'��J�� iLIO�y��̍1`�v@����΄!�����Z��B���"Ǜd`cu�tX��K�b{�FH�uu�~@���,��������W}�C��_c��/0S9������G��:$}���1;g����v��jD>8��.�9v(�_�������h\���FӚ�~�aD������F�FI(�V-�h�J��K�V�B�SW0%�xɋ�͈̠��' x�(����8�sQ��`5�%�ڹ��B�*4��<K�Z�?�j���\�G 1Z�/4g;��`�H��[J�$��:4<�ȃ���J:��,�.���+�~N+��F���4�D�� �mw ���]�k�q\�)x��drɧ��&/î`���+�:��fw��,�qt���m���B�"�Z��i�[<�‵�F��A;)�xB����vGzbAto��0򕦿����>=�;�������u#68��3���U���O��%���W�s��N�	�V7�h����������Ú��� iE��W�F#�]���]C�at���t���n����u���k�ι�'�玔�DV�;Q-T��K��=dԋ�������;��,��hd��?�7�H���ZmM�G��a���e���͔��G�(�4�|�n;����fճ%�q,�G�����u-�� H	T��Qd����S�����Ӹl�-W�^!�i��������`��m�pE��@F���'�P����Gp9�)�l��?S��cUךd1Txw����Sl�&��z�!�l��F�d��GD�&ӑ�'��ܟ߬������p���o��1;�,f�6=�C�~�/שOat�&��[^���Z�}������4C����.Gce���G%D�;bv8���6�����H��̪~���"��?���z�[���M6yYAq��d��d/;;�q�Og�vꏬE����m�$���Okى�X�]�<.�!uҹ��\���=H��8��)1zv�-��+p�^~m[�|Iȶ1_���k�9D�~E��zߩ�L�!^�OW�)��ѓ���B�<r����{Z���q�˭2oKC-���#���������E��^ؙ*�Y��Y!��~%k�����s�Bb��Y^D Y�8��e�nS�m�&D@`%�'d��:;��?�Vς���>�;�K%.Tط�m���]�c���sl_���-vto���h��Ai��d��G��]��~�}��˼��HF 3����.PJZ�����(�W�,�9왡b��'U�ɡO[,�S�汝�@/"�Ӿ�Rs��n��奤��z2���Y��A
�e	��1M&�4�_A���L?G8R���]U̯(��e����D�L:{$���4n��Of%���J�����`�5�C��Ys���^"��ޫ��x�V�R�0D�J�&�ҽ����vz��d��@����Q3/����Q�'Y˂���~�H�b7���8�pZMt(d�]=j���/**��	]�kQ:R9
�U�'�m~����TtGz�"�B=�6$Z'���M��v���M�Sc9�p������I,x�W��L����ȝ!�=M��S>�}�!g E����)�]�M��ג]$��)*��B�7��UfH>k��`&�f��]w�t������p�\]���C٤]k�6P��lݰl?�O���n�>YmS?�_l%h(����l��7��i�Y��N_����w�k���Ɗ�t��2��X>����o����z���cY��)I+��c+���Y<���|��XJ�	���bn@�e����U�7�9gd�rT�ɻ����漎h�|��q8w�p��F�e�rc��	�ǭ�P�!�k}�B��I������J��i����JS%D2�#b�q��:9��:ߍ3Xv!���	�[iP�mY`�L�2��g6��\:�� ����HF������O׋��IO�`e;2Y�S:�.S���>~��ֵ#&��~���I���ir;h��=�g�2_����S����\��͓�������k&��:������a���6�P[�>1WZ��9��gB�3-+��=J��CQYy����fBB���u�\��WچG��Q���]r��=��D��YG�}�4�s"SD�t��	K_,��I_���;e�a��wБF�w]@@Y
=�#<[�fd�خi�O���3�};Wi��;=��_ĭBl!���X>/�N�������������P�S�1ۊ�$��Wb��Ӯ�t:���Q���\�WJd��%A:#�R��³BC�eA�6��GLJ��#IWE���N7IF���N����bI�W_�\�X��������͗dkv0Sʁ������T�}uQӈvUM\E�)�g�*��j�V�¤j$ص��ә��F2�����p���w=��rg��:��t��":J"W�i�>N9�j��~>��v��_7Be���џ�������l�� �h3I���Z���
������%* �I\��x��y��Ѝ߯�n�eiQ�8�_��e�]������-�Uz���P.J��c����P����A2�#��w�l������M�����W,��qq�c'����+6#75�i��8H�u����>)t�L,+^�QA�HT�+r��Go�X���a�������6ۇ\�ȹ�QRE��Mv���A�z&mN�
����=n\~e,����݉�bx�h!�Me']�����O����5Ь�����Xi�
󃞬[�L�D�����&��8B	Q5�?PP�py���յ%��ѱr�X	m�vO[/"��kQP��iĉ�нy��k�ڞ�ʿ�`��JF��<��$9�ٛT��F�D�B	�ٔ&�	?���aS�-�ᩑL�!�1��eJo�4�'i^�%���a`-م�x�H�Ub�!���ڗԥ<`/��U�@E᧚	�p�}���gi�"\��ѕ{O����2��a���J����9�M�r��Q���6�˰���/4@zG������?���]F}�(��i{H$�%D��'q�k�=��nru0�{�`:?*�ip��jG��¢{���X�O��j:�r��.�GV��og�n�^�)�+�!!1	��=N<@OA�z�y|��@��R`ӭM�ǻG!������iq����3Υ�BD����m�|?1B���K ��)��U�k��3$��
��#٠Fm��yO�˖
$�	rU|b�v��c\�y���Ⱦ&�"muKGU~.j�^���8;����f�Ad�?]N�ߒБV#�.+{�H
re㵡+O���b�'�U�e�P���l�*0]wR��>L��(:��a�|a���e��{��������GsMMgG?�#���J�j�����'ߕ��P��q$���T�8d�J��%���=]r���ԕ���j�_�l�����^�C�~����	�̲ZM}6�5�Yn��U&&3[wXp�gT�[��Ywt�������$P��B���vK|
T�����P��ͼ]<]�^���~v;k?�l��'ik�P�)��V:�ƦSm>, OUVv�Q�s�1��iLd��P,�A1>�'y�ᦵS��v��K}9���o��Ip�Z�4��a#�DYPF �.��<����Q���
Z�^֝!8�w���I���#e��[rb��#�	)�E&jmH�v�/7��೐��s�E����	���dpG�T��s�=)�~�O����622r����xmT�V��K�x�����Y�`0��jpx�8�O6��*]žv�ah�Mխ1�߭	]�X��������4��jր�,��M=���?ټ���S�L++\�8X7��<�[���r���x��e[�,Sw�z[v��`��o���;UQ/�M����$M�&��a_v�b4�g���y��1����2��|u.*3MUg�Mq�Z�im�\�H�,�{+���y��)X��zU�Ĩ)*�Du�n�`D�$�ZW����맠�����n�>�����C�SD
1gu�,�w@��_�c�Q~nwF�+/p1%������MG��_23��� #���A�R�G܏β��m��?N����ͻ��j�5�Y���I9��(H�X��A�ur_���՟�z_43-Ssr����o�dS��q�,��P�~�h�����W��î�$y�h���n��Ӯ�VE�]p˗�:o���b�6b�	�:��4�jt�N�\p�8�C��\� ҡ��|��`&�b�S�}������ƍ&}�ǉش�>U��;�����Uj�-��5wx=e�Q싅��JˤT�n����[=�G���������v�7	�����_{�ߤq��]�N�� �:���K$4{�ufHI�ec���.�*���R�	�������T��Za7���y�y� =C�_t9�ڀ2�8����(��p�w�Rp\�z�0�-��M�]\Dp�}8�+��:o��6��N�e/x��H_���
���v���h
��5���5�ǋg�Ғ��o3�L2��|���|6�Nܛ]lfJ�N!T���-.��Jk��+E-�q�O�d>�Ă�+���OBսsj���߅	+^��s��-��W����t=ed�s���+��`�Xliƥ�n:�c`̭"{!�z���M����p��ŀj4��B�%����}&��nT�
n =���Jm������n���L��Ԃ�~�� 
w��&{�8��'����]+2�G��A�6װ�ΩZ��Rёp���|�B�<�V��$���ȸ�z>)z���L!nJ]�NB�p�D�����>��3ˎ�lĴVavƸ��a�Q-�W&[v���-�PWSs%v������o�?�����)��|�K���m�OŘ!Ҧ��1�X��҂��K��_2��05�㳁���49�f�J�O�����g/��2y�J�3P��I�*)�˻���׺��*���-y���Њ�?���v�g�;�N�O��>ݾq��KJ�W;�ީ�³��<c����ޥY�!���)T�g���ړ,�>
��7��|T�AH���������&G���LDc��I��NM##�%i�}3l�R�ߴN�~]c4�V2>W˂�A�P��w���6��2���"�&��.B�ml�CLd�"1���b&����Q}�`d�\h��_#� ��Hc�͔��$���:�M��4B���I��y�I�j��V=�/�<�w�DC�9Z�ppww�JQ�n�
����)
͏�����C���@Q��|i�"�^و�3�h3d�B٣��dv9W�.�.���jbb������Y��{)N����ŋ��
#C}��i����v���14�gf���Ṕ�lyq� r��9�ɲ7[�*��߅&���si�o�M���������P�Y�Z�×~v*��p΄�ﰞǲ�U�ͪ�$�{��h����/�ӂ ��.pA��:��!˞,�%�~������X��i!V������u�v����M4�9(sVe+�&�X�ږ�56��v��/1�TK�e�xD i�����9+1+�����	7�B���)�~9[�= M���S�8H����<��-�E�fw�.?3��n �M�!R��Q���SYp!Ft�/��6�Q�X��ֹ]�~"\���Ek�.�Z��PJ����^d(�������<�x�1�y�����g�����,�	<|�=�|x��͊���v�C�����I���k�-���fv�&�W%��q'�=��[鲋�����H���($Źm7�_�v�h��;�zZgG����D"k��?k�8&]'�u�DD!�M��@�V,��G�&{Q�J{~�8�����.��X��` ��l���b2ƅNߵ���� 	�i�z���WBY�u���Ѣ�	��Y.�ڥ����G�'�Ȝ[�h��vU#���橳�I�J�� ]r�m;���X	Tt���e7���ۚ�r�tܳ���]�.�Ҥ7�դ'�������͝����k{4���~i�D�q"Y-����D6x��p�^�F���/���T�Qs��>Bct�՗�
��˽�_�,$Ex�3Ф}���������~�K1>Ue�T��'�cXl��J�,���Yca�LZ���U�H��P��]nr{��N�`��n\d�ZjГ�SȝJU x�^�Yz.Լ����k����g-:n.��C�0P*��#������f!j�G�2
1�'�b���9���d�{��%h�������/{�Z[[�@Z�n��P9�*�tE</�R��&iV�xL���>��diZ��wPQ|�=��9I�'��q��➿�W��_P�Lb_g�2d�ퟷ�Zv��;Xdn|�?���T|پ�#�V�XRH~M�sY���ґ&��p�5�z[�TZ����-H$��;&�B�W���/9YM����qm,�r�t��ӭ����'��0��R���I<��Yn���R��RA���Uqi!�L�ᅛ�O�N��%�ۜ�����X�����yg�y����ʖ>�t+�YN-�@d�֩W��<���&d�HF"����2��ط��o���[]a�����!�����
Vx_/7���j�6�#��@	���BN�E%4�(�y;;Y����~��'�$5�\�c�&�o�k�R`��2�_�/�u8�TN<�g`��MkY4��;7���%yz�!WZq���U��;������b�FB��O����:T�}qќ�X
C{�C$��HZ��=4�Yw>�ٍ���&�S��f�J�0��rS(�ߌ���C�[����������Z�3���5B�K�ѵ�p�����O.��-2S������s���|fѩ��[j �ݴ���Qg��u��Tߨ��;܉����O(W=� ���
r���\h:�9F~w2��`�}�����_���4�������XZZkí��}~8!'e7�����%����vW�t����`7��[�H�� �M����1|+�%@e�l)r���� ��X���.�P����jc���ʮ�3�,BB�Ts*U����5zo����YEA��_6�;P��z�GRS�G�;�7�'��р@����!W�zyM�'1�J\0��ϥ6�����CȒ��5\,�ط�.�<�����'��&��.�������
�[��S��8��䰄t}�V�%h�4r}ğN�b ������OY~�F�V�y]���^����^j�r����H�%����1����[�nOp R�[El�&6JPD�,Q)�+��{�}c��`�=���%���xY#�s]��n�J��[��\�a��\ݚJw��+���!.d,$��F��<u�5�{ț�*�k0�Z߾I��T3��G޲� r�v��F��8�@���Z��Z���ڦ�%�:f~^\\a�v��D���1ª��7����jn@c�b|u{���~�Cvo��ǌ��'��J��L<t��տ�8�OJ���+�b�q�W?X�_������ ��TN.b���vJ��V����,H���I~ٛf���K�|��B��x=��t��!W�y�~����c�����~���̝�d�� ֭��(_�Ɇ��7IF�t�XmU�-Ƙ򒳋KR$	�q���}I�V�����{�UCV˰���S��0��M��S����Y7��-�9�{���sۯ��U�G����S��r��-��[�������j��欹�o�WS������fv1���jˊ�(�j�f�i���E��]!���'1�l�\�������I�Vy�����q��A��� >��� ��^�O��n���l���$@_�����b��v	�b�lD�-��?T�GX�J��:YF������lƨ������ȀC[����C�I�H�]����<&��<®�����=��������+o�����?�J�.b&~�b>�H���a$=���r�b+C��;�Pu����O�H�Wp�1��ȴ�P{���r5���
R�g{i�ˎ�B����H$򘟱1q�ֆq=l3���у
#�2W������� "�m0�NZ[��+/�'L���M�8N�E��@r��<���� PHf�Q��y��b(���Kv|�`�������&GC��&�YY8ɇ�xxZ��v���<�;�_�y�H%�p��G����=���r�U�����t�V�����ng4�#���f����B9w�[��Ëqw��G&m56�K�/�b{���kH.��#�Xtɓ6}n�ޟ4k&��K��Us��R��dX�N.�<�س	c3�HvO�ʯ�'d00,>Gjc	ä�@��"����R��A��k����.E�@�dD�:��;�j�j)��.��9�����8�ɥv �	�ju�"A�콱�	���U8E�������Q����/�F6����9��[]�?���*��$����1���R%�N�Vl�6,� nw�_��k1ctK��%�T;RV���|m���k#��(�H�>�`�ͧQ�t0�{�μ�v�_��Bu���3j�.���1b}'���1j�g��3]�uQxS+G҆�������г{���E� ]{~�
��r�48q�4�N(n�j�
3L�`�M��]�蜅?�6����D&�Цz�Z�sss}��F�.+U4;�Y{z}G>��*�>���q{�b������_ ���>pީ��M3V�V t�\������먂���60R4��&�rƚ?KFA[t���O���&˅��U�_^���2�L�m��]��"���|w��Y�e�����2U	Swz־^�$=م�����YB~QĽ&tG�.J� �u�k�I gs/�OIG�t�݇O�
�B|M���(���5D�p� :+���'@s�t�]�r4;榰���k�7�����}F�Ff ǻ������E��^&�Wn �o�d�;�%P�� �鵛��_����%`��L���M�7�3�:���ǬH����� 2	�'���U+?�(Xd�W�f�ə���
]vF�.�y8��E���H�_<,��Mdi���~!0�+%�!�l�H�ʋξ�w+��$O�u��̆^���bvB���+��v�l�V�^R�@��r��^m��9�z��B��i0nS''-J�*z��bv*q�~����;�b��G��o�78�!�B�P(Wg0ց�I�MY�I�q4���+aI�UU�E=�4{ۡ]��^�O�<���y4 ���$��;���B"��F��q�Q�L�-�.�S�|F��L�Ϭ�?DN"�&�ls�����"���%��.(�a=�>���m5�{�`�w�9ɺ�B�qOj��������~��I*��iB�v��wf�-Y�a��oϞ��.|4�G'tJ�S��qaS�L"����!�)��9}��)/�OM���/K��to0A(Zb�Z�/ʘ}:؂3�� K��hy���ǼY=-�e��'B&Ԓ y���1��T��b^���9�k���Yr���W��4qq��A*E��,�q��3�w *	�ݺ�����U������`�Q>�]ǃ�h�E�<׃f���ʙ���7��1��5Ǩ�d	Z��`l���j ���ˣlD7� ?ޒ?�I»Շ����Iq�i��d��`D4��������f��*��ѝ����,�:�� R�/�z�e	���
K�;j� 
\>Af���o��8庍���*��{
E9y�R\�}*u�'�90�D�D,+v�1䔌��N��r�T����L��F����	���k0x9>��8���"��3O԰�r\�|�3�J������.P1	Y+��+{��Sط���%.�E���$V��������Vȩ6�B�I33�~�\�0�R�
l�\�#�8��T!�nv�E�찳�A�ǁ�˳O����prjV����_��Ӧ�Cb��"��,�S���8��`���J����O�����t�K����Z�f�.
�s��O;O������D~�F�F`7�d�o���?���7P���A�|R��o�!'��������>987M���hV�G"��w8���T�V/�Q�`�c���d.��D�U��ز|��<<<4bN4=3��9`\p�+�(Sb�����TiB�NG�	.GRS�6��d�E~o!;��%'Z���9���(�3f�~=D��#/;�!X$�`���;\�¼���l��k�FaM���*NґHD	%�6������b���>\w��~��-秱\�h��r�onT@[�pm�D��� ���B�9�r<�jLR��f���"��f��0���{-b��(`9�CHj�eT�����#��F�I̐bM�1���U�{���=�y�>b��ܩ�~�X}�����	NX���j�O���������mM�J����*,��a	���O�%���ѝE�br�Z�I�X���oT����G���/M�g=%�_þ����רE�yp�|*O:n"�k{/I���G�Cu���:	}�u��G~>��.��[��r�� �C�q,�V0JU�=0L"W�u�{!�l� 6~Y�q��h�d�D8�%�xK� f��Z�G�ѕ�Z��T���sTQ}Fy�s����1����NZ��/)��GTw݂d��8�ő�����%��V^�����r)��a�����~���%�����1��0
`�#ݨ8ş	I���^��n�=��\����<fj2���~O���
�\tKxGBp0ɝ��ؕ��4��&�����x���Eܫ���w���T��¥X�Xf�f$]����j٥M�k���>�#e���p���yMz"t�]w+\��^^ �;���͘r�QǈHR�(ݺ��N��ջ+]����S{�G0B!g�Y�]�p{�=�ǀr�t� ֏^`z�)KRO++2��� ��WA����i$�~�4�fH�5Ju�3k܏�Y���}]��u���]IbM�^:_,p�������{�}�f;�1��0:H'uZ��8���a�%�np����7�8���'U�����_��(~�������}]�l�Ӝ4HS��G���ǐ������RuT>pXX�K�D7�/|�)��5ކ���a�����=����=ky�w��� �"7��j ӫ����XD����qH���x�x�ɧ�;+�섽S�Q��f
R�}/c�H��y��&���{ntn��q�W27�\Γ'^�kA=+o�-�H��z�_�S��>��S���5�T���H�ؔ��@p~�F��;a}��
Q�hJ����lu���$�,��d1HF��hMҎ|G4�|��Du5��:����e���AC���
\&FX��|��������~�n����2g0���'&��z�%��T�����A$��&8O9W�e��n_6�9�'H)�C/��)����+��6���<��0����O9/Kʷ6b|�A&F�[���;ڬf��=��W|&a�&U�.I��@L��t޳Lx�12��T���F&Ϫ�ޅa����P�{g���}	��\qE�;ݥ����CM��-3��4K�k.�,��] 췥�a0k��-QL~�n�^_�DЋ�$�qW%\X�5��@�!��� 6÷�t	�SE���Z�
>O�s*�!t�P�o7XVX��[�Z@����t9I��(x�g�H%���������ր ���E� ��$�4�^��-ԓ�Ԟ��,9�&���㏢M�"��"�Ens�J:��^+Z�$�۰�U��	VHgs��ĳ�Нi
u���$�o:4��ï �\��F����B��Ae�c��h ����_��s�5�ؔ�~��;q��sL��U��=�?��r��.�����Rl;�5����m��j͖4�[�!�Q� a1�	���"������<�m(y�'��u��.]��P���D�k�~�	]q8xd}ϩp����Z� �@�Y٧hm`;eWD��R�p�jr=z	�̵X���:k �oa����_������P�Z���n��rg���}G��u��]N����r,;���j�������c`�������w&ڦeM��*�,.��k�f"��/΍�'Y����4����.���
��� g��|T�O����ڗzዡIr̐N�33�$?*�����x�>Z_&������|u��n V��N�D~)��eZ|�ZL|<���o�B=��:-�Wd�->y���kƸ�ҹ[< R�O+i�;  ���O�W|f\�QS�\_F �f?�(+�;ٷ�������5�珅l»4�l�*�?�-�,*�dd:l���O�;#g6ۼ�c����-��V%3���s�x�l��EK
�6�g0�xN&���4.�ןpi4�6�[�+�E�w�<�ϭ'�S>�k ��i^)\�TD88����P/\�anT�>��1 �B��{Z �K�v<�]ȔU�riBpW,��Ȁ(/^	������%��pj��{��Ŝt�;��ژ/��oڀ��#B��*��k���� �؟�k�����;?mD��Q{����R��4çE!��i��e�ߞ�Q����ދ��b�"����@w����%k�wY"���z]t�%V�܈��j��$�GNj�X����a�eE�	)h/?�M�,�&�Рk�k4��0k(d�q!�8�SzӇ�I�A��U��
��b� �~��s�U��P^х��V��O�c�a�,����M�"��{��v��x�3ԫ��U�	�k�����,�kVX���hMg�m1�P7�9�&d�A�l����>�; /��P��o�M����-B���������������x�,�ʯ2�R�SӔ1Py��������E���8@+����^��fw�����Z}'+��go"��U�aH5�sFm�4O��{��ׅ"c��I?+.1ӸF̦��6ȆI^)r�/�������#���Y򕯚���<��u�G&6+���\��\�f�K�����FOU *�𯳳ʗ�[V�\R��	����	u��JnG_�Ǐ"�/���/ϼ��xM;�k�m"oW���]����V� �1���Rެ=�9�%���pP�  W��W�Ӗ���T��>u��%�.�VCsu���yzΥd�d�N$I̵r4W	c
�8����s��&���-�#�6a�{U��w;�ɜ|�!���ج�f�;sp�ߦ6��]�T�$s \
͎�����)-z��y!{�mvmm:��`^,�������j1=�����e�Y0�g�:g�2sZ=	XLE���] ��H�1D�0&�rA���s졋�QaG}e�,���xN�!^!W�����0l��Jmnß��qĲ	I{�H���h��Hͳ~ 0��֢����ݕhVV!�y9���Ց^�����éa �j�;ۍ Q)ҠR�M�s7���Vd�n8�e�q5��C�
���KJ岱��.z'�7�f`���~�3W�7�Фf��G��+a��7��䭜�E���/��#e->�O7�������ʃ�J�z �6彔R6�Wx��uy�]U����&�ҽ�ض��%�Љ+H+���H���*�� 5����s�l0�'f��L'j�����hW��|@1������?�X.6��hPُc�-3���e�WMó���e��)���;���V%�f�jz�m\<�!g�͸�ckõ��梭oU��x��+�����7���>�J� "��h6_ek�w��s�'��9�����B6`�Q�͇'�5ҔS����|�V�����;�HS;����V{����5$^�,Nw�b��G��>����W}}AE���x��W@p�V���?s�4��������+[��V���N�Zd� �������#8���̲�v��P�i?����^A��K�#�/o �I�`l͡��qs+�3u�<e�I�sބ�g�i�L�w Bq�(���Y�����o��.ZZ<&!����Q`���ӄ�	D�iN
��ǭ��5t���?�Ȕ��&Q_/?��c� ��MH���?bz��Ý1p�6
�O�3��`�j39�(y. ����H���N=/*0i��s�=��ro�B�.�b��;����_'��7�,������hi���u�ވ�A'&#3R:I�0�4J���	O�GV�x,^�H��ܻ���������v�-+p���w�\���!��3'`y˙�7��$��Y�IU� �$5����U8�V��ã;ö���6�y�sv�_�|>NQ��EҀ�F������7��d|����BO�L.8�A�j�e\B"�~_�
���Գ7H� e_@H3��bq������e��PE,���_�s�w����h����9,�]�2ҫ0�nF����O0sI�dd�|�#����}�n�#���
����bk��f��3�x���Z0��'"4wà�~�5:T� Z���#[���rߧ���y`??(xw����_'�n�v�w-���+4N9܏P�w�.��#!)?l)����f���i�P���?0*k:3�Nf%,`?9;��6� �k��G�vQ�I�``�.��G#((��z�/ϳ�Ya��*c�Vg5�=�E��ּ�ۗ'��.��%�cErk
-�j��9���3��=x̠��p�U��urEL�Q�;n�ZXu���HO��=�0jH��8N��攪I�n���9�_5 �{ڨ��:�~��^�C���u�S���
�b	y�^�J����e����*�S׾���&�d��_^�����B�g]��:�F�+ ����Yj��8'�?\^����6e&���(�m֮�y����'8����轪�	Sg�Q�ww�w'�4�|=!d&1ҟ�\ý��G߽��u8�Ô��sak5����._�+���o�Q_6a�N��==�Meȷq�M��������ϣ~3��Zn��wգ:"�_Pע��5�%�9px(��k��eF�κ�7[X��)�֤rDǢ���`]i�S�!�o�:���}�1N0��u��9�nS7�ҫ�� �B6�G��H<Ę�?ϵ��*NL���^��n����^���%������������EV�ɧ^mEi�U����1�8f
�����ce#��F�n�����s�����ځ�Z��FV����~t���� �dM�"�'�:�y���-�mm��\/��&2���)�`�
o:)���n��&�_� e����s��g�#&��f���q���.�
.�vn�p�7gy��b�|�+;Q6�*e/)�2����(�Ze2{2[��=��Y�R�P[Ż��dL��S��C� E0��	��T#ʃ]�I-O��uK�@�`B���y��Q���dx��/�;���jɪ��[ʢ.#ܼg�g�\���q�S�}�2I�^���J$hP�L��P�S_	W5!>UY������BئExȖ�z�.�,���m����'ש�=T�6vz����\2Lnc٢���e��b >n�i}�:I���-���8�+)��C�B��ʉ/��je���ާD�����LM��ln�����XhĹ����?�o��KGP�V���`����h!����I�����7	͑�uFZ皨�j�X��롩ȶ����->7�X�����N�cP��Yԅڥ�q���y�	1�/�I�.b%�����
2޹��#��j���2����V�}�Y ��.OV|@C�ÀW$(�S\FLǘ;�S0g�+������_u1����	PlKA��ɱq�G�~}������ߟ���\I>����[��}���Ó۞�3�� i9�Ͱ�q�_h�I.4-�F�] �1@.:�_� ��	�΁p��G|��ܻ�d��У;X���Շ~���)�ΰ��� �*Ǭ>�A�9b'��������)��h�J���O#N`�N���%x)1h{^��I"���,��^|�@�->�(����Lx����n�,_gˇ�#y�3X�,���KJJ��㲾��_��ҧ >\����V���?"FR�K��Չ	�V+��eN"$1�?�>E_��9�Ջrp��'h�{�h�f,��E$&	���G4h>]�j���#�ڤ�����#��	$���OH�}j���P�@Oܼk�ˆ,�Y�4p���F��vb�V��m	�_M�L�l&�z�������̂?�r<���չ�����9V�C[�+�]�3n�y���j\�ƨM˔}3�,�i�Qb6��c�P�2�\��.��
��� ����^�s���Y�"���z�A���I���8�cT�e
nR��L���O�؋��_z��~U� H��H��G�����t���8���{��>�QZ�8��a����裧tr�)M�E)Ït�zl�dM�I�LKMm:�g9���)�w��<[���K�7PߞV�{W�u�QgO��	`��܊xG�%�΋x)�.���[<�~��M�)�z��i���V���v�!���p�r
�({�^�3+��S.|�p��G���S];�L�5�Զl�T�mc�
(@v^QY��E�{��.-T>����߿G]C��ɨ3x5
:�[���z�N����6�X�h�����l���+�z��O�Y^T�^s���~+%�����m{�%j�u�h�7���%�1;�%He�NHu��2��5��ʑ!N�����DolR!j�PmM
g�O?u������緳���m�v�N�˕�l����7�sT���K�dznL��3ԍ�JU�� �S�f�l�ړ������62�6x����`�d��&��$e�*!���t=D�;��|�^^�{	B;w�TK/�_h�A��1��\{i������62��+vdѽIi6��\�F�F�ǏXɲ2���~B��js=A�;�f�����x �5Ie��&[Ti"��$[��	�+������V-�w��uX��j�=7�ps��^��|����	1���R�v-�\B\�a_�5 {^aϏ$���%�"+K}�lcƚA��Q�T�p�!���M�;��9]-��M�A�{U����	Y�^�� �����#��nl;�ض�_vc'll۶�d��7�m۶m'��_�~���Tj�>}��ӷo_*z�vn���&���x���#������شf_L�s��
\�Fu�����8�u&��FXGvT��@X�r��E�T)�8�U�+\���*9��T%'g�����8̀7��o���T�6���FL���u�%�M�鑑�G3p�[	,fCi����AF�^��p����-���]���x Ƚh�:
d�����4�S@Q�7�e�%�TL)^�s��V����pY������w��/�qn�J�A��6��	�sĖ������کF��	�΄�^�)7�\}fh_ނ%��7�!-*����ob���D��Y���;�8�F�b���,�����o��W�_[u@�,Y?�.*++�+%�^����Lx0�����Ow��*�ljp�Zò�yҨ�N:��vl���z4,���%���a���n�r)�=�QjI���?��6�� �_�!�:�Zj�Sg:U�x��wTTX���/MT{�я.Gb�>N�;3>��q�p�� U�W�i�'2�h|$�_�n�M��P���"씵�Z� ������b�@�7������v ��㹹�Ab��l��\Dd�Z�$�^�M����հg���OIA&�3uW�ES�2z�
z�0�+#�(y+mF��5�w�Junj�|$�R��%%%φ/=�{/֞��t�
���c�I'��Z�KCy��bd�R��΂�8	8�7YF>�?����s��;F��B�BΧe\���V�6ٽ��9�E����.���T�+yD-~���|�wm����U]|�����J���{֓��O�5u⁝�~���X�d��U��l��PD��s�u��Śk�ԑ%�C9�!���9ϳ}L�}Tg�F����Yۿf��(n��Cv�X}����M�����@�155mí3���vkg���xӭ��.4��V`����3$�Mu���<��{~'�8�?�^�� %"piعNw�",c�y,�	�˩]~����O�p�]�|i���Q�l�[���r)E"²]Q�N�� ��;R-6�w�k�AC�A�Q��Xk˓������(\S�6%��aESSs��P*��5b�8J���6@���|�� �;A?�N�n�Ɋۯ{��z�A~��u�1CŹ����|��Wȣ�����U�r� t���eKW]_��ɴ�x����@g�7O��,�@���]`��5e�>ʶ�|-��B���ejUlG�YoJ�8��z�7� l:ވ�y����� �L�1��PN ��5#�L�~1.�%S  ��lP��P�m����攫�$1��u�|�iRu���� o�Z�56}����ҵ������lQ���ܥ�n{��C��2|W�0�����!)��M�lr�G����˱�	�p+曳ς�������?CD���g1�!/4����_�l�i_OM�_�w����s��{q���}y���Oy�ڱ��������4`Uu6\x�y�n$T��q$������=�oN�/Z�F��a��=Tu
�4����ǩ��h���K��Gl:�iL�~���A��F+�����c
7�9P��H� j+�i���yT4I[�������-y�a�!,na��%�$Z��ޞ��U%z��o��J>k�
��3�F��E���K0�x] m%�s�/ ���������η���%N���/ӡ��,�^�?@���9j��f���TLy�b����1cZ�C�>����*uҺ���$$���T�03j�Y�Zuj��z<�����~ݓ�5V��, ��-�-Rj��0�yXԴ%-�)u3�tſ����
��(A�] �W��x �ҙ Pia�ޟ�%J�uf����J7�r���ꥩݢm�$7h�~4RPQ��O�"Go�5�d�`����M�n\�ޖHk30y��H�(��
�O3�!S���*�܃K��d�^'3�TFr3�W�e�jgfq���)b��R+���߉�שׂ���^���&@p��f���7���
��+�,J�A[2�����d�ZA�$�Ew��Ncp�JP��B�W�G\8)��5�<S����T�Ѳ7޶�%�v��^ Pc��d9z�q$�0^�d�T�W>�� 0q���Q�r�A�mg:�ղ�\��1���D&(/������l>i� �^�����8۔�t�lFO���X������m���䉒��J04������4H�h�򼼼�=��8�$<�c�γ��� +z��4��&ǩ]A Vb�$SN��~H �h�3P[�Y��vD9���a0!�At�)T��,�������q�7�~��>��*�𕸰�_f����u�p^HKMmz���m�\�d���](]�E�Ê���sB�#���з�r�Qj�A����'$]��3�U�n	��:��kŁ\��Ԭ�Y^�@��)�H�{e��Փe��qYv��#�@*���]RLM�V
���l�V��a����_Qf*y8��	�k{�b�$�2����?��Q���T��V��g��[�����_�4j�R�z��\����!�����Ӭ3W�嫵&۪����K� *���*��*n=-��m�%R���); `k� ��v���-�r�G0;
̚�Б�z�p��r�DG�����\>�!��_�����~���h��Q�Uj�8�V�J39�Ida��*�m���㊩'0��>�T�����J��eHM�X���DE�R��}�i���Ԧ�9�p��\�T.�xp���jiFlQ������z�TX�^*p܎�/��}��}d��0$���K³�ۨ��#�d�k\�:+U���ԴJMA���Eb��E���L�_\�5=�ZVM�n�C�� �3 ���@�Ļ@��9����PZ�����+��y���m��Ne�����~ߠh9��#�nE���i��%G�r=&��PB��VӠ�y��X��4�
�!b��H����t���l�w�ۍ��1�$��؟�W9�ǀ㘢l�o�[�h�V����f����K��*
����ᴴ�C
"�
Y���\�u�c/��ui>����*|0&>��i�c�$3������7��W�g����dZyO���.��̇.�;*F9����-^��{ו�y�GD��'�z�n��& |�\��8� ����F%Kz��5�DJ�|�XY �^t���$弔'�mi� ϲ��@v��@���A�8Q��M���y�X�(G%Ð��mX=���kY��:�^71�����eە�tޟ-��0Gpa!����RK��;@7�c_�Q1�;��j���Z��8��5��`�8��v�=�$���BX�"��*ª��mJ1"<��w�x%�,F.1l���9�b��ǫ	��^��Ld�8}u��W�J��h��ק��4	��O���G!S�N�i�4y"Ml������7�i^b�'����g4|��hx)�G�e��Ȓ�@ z��\��'����~o Q+6�l���ws�LAR��(���Rp���x/�(�@w�	�!���7JNOoa��0ޙ���o�^�]�?��\�wm�h0����z=-(HJ�گ��l(���\�Jl�}����d
	���T牊����P�*����4�}6�W�aͻnf#|�6�n����4��ĥ��T��L�14n�l�uO��A?.���+���iH�(0�JC���4�0MS��D���C2��[����C����G�M&D����pI�@���(ռ�-s>[�"��9P_Q��uc2�O���rs��/^b����|.��D^���9�.@#4���G�n0��Ȍ#ɬ�� �{���o�?U�o��0�Gm��u#<S{��U�͒�����V��*7~�r��1Q7m�C˚�S���h=��8xr�An�KՒ�j���F�Zc8�/��Gi9*�~�x�%��)�Ԙ>�		*`��!TG|� ��TH'�R�Ǳ��~�@�:�*���l$��^e��O�Q�1���AΧ��ZJ��1��Jg���*T5�!D;[C����6�}w���u��S��/9M(�㾵e`�[���`A�ޠ�@��KV�1~$6''t����� �H쭯�����>�Y[�zZ:9���C�����K�Bj
�@�ЯU����Co��S��p�C�026����,7�ۊ��B%�R!����W�*H�ZE��Fs�4����dp�;�!��Hz�����|���N��!�B�ȶ�((�a���A�b��� ����_�4�/9 O�h��֗�䭟��A��P�z?���$�>��B��?���y�lm ��>N������x������`�������g��o����wY����x�P���lI"&�8�����;<[ , �����P��Թ��9���aq��>mLZ	�i�b��\�"o�?�nhj�S�X�S�$�#�n�9�'�w����Z9}�\��M������-/����`tg���\�>Z9�\7���<���AdU&s~�@���$��y:�EO�<��k:��Y6
�7�԰���[}��ٸ��K�#n�o�*3낗�7S�H�[�����D}²���x��{*�g��b�&[���t�FF\dA�C��_/�����i#.K.G|ݯ>��C��v! c���u�g37�[ˀF��=vhNïǌ�63�(��$��`����(7��)�3�\u�5* �@e�$$��PP�+�_���M.'�R�����q�*K�ͷ���~+-lz�|9�����g���10���׎u~��2j���qk)�����u�UwS_�	t�\�:(�Ճv߬�<g �j:-Ue�>0������_�O���M�v�ec����8*�}�D���wjbV��@`+�e�����}���F4��E�V4��C�d�``#y��B��������s�৩Ѯ���m���������<ժ�¶D�w-m���j�b��^-��-]��$n��!��P~4*h^ZG�)�ȡ��*Պ��]:�x�����M�=�j����i�A�o��܇��̂��HiA7�M-�u������V�������ZSBff{�~_����|���WM[-�6i�c;1��b�6�1���䮂��f�~������I�Bۈa�rA�hu��/�M��>G��Xմ�Cp������L�W�����Aʋ�ks�x���������gD=�8�M65���V�۩`aU@��/�2�_4my��[����aP7}7��h�!3�J=�^��} "�;��(�ܠ���	8�*���:���k�#*�ޮ��8��N�^��*�D?$��`^Y�#W�[�f�2��ҎlПK�Dh	���h���Z*��W�Ow��ɫz���3��5j�Mh"1��������!ړȡ�T��wtp@����,A�YͰ�f]G�����t;a��$%9O�vߤg�G�	����0���bS�M�\�c?!6���S����+����_��^�C;q�1szBl:�*�A`7��[�m�"0�B��θ�]{]|�2a�S�9ե^���r&_|�N�����@��n(������\/ػĘ�����H ���0Yl��0�m�9>�
[	��7��1?��%�K]��J�h�#i���9�c�#���ggə�$;k?��V[�5MWj�M*@8��%;j�h]v�A�p���h�MD����v��Kꕠ0��6:Y�����C" <QP(�����g��ܩ@�\�#"M�?nI���D���<`���3�\(U���&K��㈊�EpT�i���]�}�����Ri�����ہ� OL� +��-����d&|�:�N�s���� ��;�LL0�q�/o3ۭ�:.^|/�a�~4<���%��e�!��݅hP���i�"E�Ps��l�7�bap��I���:�J�C����pI�~fQ	���vr8<�Z5-,��X���B��|\9Z�z�ݴ����J�3�b����� x���:{q{Wm�LLL��K�F'��P|�|�щ���T��@	�����M�����ߍ�"�V�Ő��QS�h���8⵽5�b`�lF=�z����+׸�<��$� �ȸ�a�S9S��Q��Г�T�c����`|V�S�$ad)u�7�ϤX\�	�
d�=�5&�.l�o��n%C�_�.���L���TTkciz�!�����{���qJhQ�Er!��f/�$.������;���j��+@`�a�R8}8�cB�t<,�Tu<��Zq�)(FXb�p@��Ԩ�X=3�6�.��v�'{��>�^J0d�����x�i�C��]���j}V���������8�q�vo�c�����N]�si�𴱬$��8��5�ٕ �0�m��ܒ���UBܾ7ycŜ�!���I�-l,,��p���Y�Y�&v����3�l.ENT�q-Vi�1,�|z�g��F��{��E}^v�U�B��Uͧ?�ŤV��Ud�V��!ƙM�����+�I	���T�%��qRwS��e3���_�.Xm�}I;�}���y���v4w��=:�5Z��8DrP�j;���*0�� }��(L��v!�Qh~�b�j>��B%�v�	Ʀ�Q�{S�Q�֡��\#rL�=���Bs�R?�Mz���|Rc޺�T���OB+����V
,3Np��Q��ښ��֞�l1'~�w���D�$}WI�(<ȍ>�D28���""��#��x���V�&���0�����<& Һ(a6�b]�3�bUbof�z���R��kԨ-Ζ��t�ֹvB#�n��\�H�Bg�'P;�	�g�a�?��ÝU`�F(���mi��t�?Ɔ�8ό̂�w�~�A�����vq��CI��p���`!.��@�nZ_X[���=�n��e���R�x5�n������͜=�ބv5�g������,������؝��;m�p�i�p�/�/�J�;�f�n#W]��>�,֯����+�W��J��4!z=y�I |���fn(�j�0Մ�^|/!�Q�7�|��-�!�R�>��p{�+׭V��f|?�F�%���p?�=2 0���u�Ío`5
목��Jik�2�wh����(K��sϰ����{5���j4i*Xx��eI��q��gj�ٍ�bc�|���o��kW��3%��� &t��f���!!e��zSHn؜�8k�@�<$�.D�Fۊ�x�}'g����[�Q�p}�U�Ye�<��q`O'zDD�9�F���r���P]$~�n�	⒃a���eh.c(O�%6�t���ucÝ:�����l����� (�XO��gZ��F�)��`O�7/�������M�W��t��V>17��rQђ�e�IA��D��W����c�"��^�l�e�\�2�8݌��)�~_��aR�R���S��EEfQ�3"�գ�I^�� V3^H_YP@�,����T$�lذ��V�D�&u���z���f��&Wɩi-��E߈m��W�"���2i�(0��k�s��^<<lK��^���Q���ӑSo�xK���#��n������>�p"���"8� ^{��]�F�4���)i]�'��y���&�J�7|��n����2�z�LY[j_�E���=|���w��܏�vޜמI;r����Y�=��x�T��9��/^
�F�r֐����"����+�xoh�瀦+�u�}�p2�z��	�?lx-��VNAXQ����/�U7$���cU2�D�gG(�&r�R��ՔCU ^9�+��zs�1�X�~���03�K��?Q���'B�M.tJ@吉>�K�Rnba{����?]�J�rϠ�*��r��!Է�GEQqg�Ѩ��{`�E�n ������h	^���v�)r(���L6b�g�7h��KvR��x[������T8az"r��/����k�Ը��Wo2�==/� 5�>i,��u�Z*��j�4��q����<��ut#����N�U[����_wGSLi�O�YYY��=wW�V�~��Sb��8�F�{l'�Nwc�A.|���?MLL��os>�ch��p;#�H�P��ZU8	ނ�7�+��]����)w��aXF�H��A��O�3D�]�G�J�Ws-	]>�ܛ�0D��1v4�F�E� :���(�ck��㯩r��(xF֌�@�'�g�m�*z�t3A��#�)n�Iz����ꛢ�H�Jb�Г��l7R����0��f#1ة�� $�6�:�j�w�����!4F�\p�e��l��t�*p�=�_�}<7��x$Q3L44/g���%�٭�9<��{e��-���:jAQ�4���k�)$c: Fn��T��n�IzHh��$��E��X�ScU�7�K����s���"°�]�!�A�������(!���p�6�1�^���$K�a�A._ٰ�FB�ez>�o}>&s��;Iz��CN��~���ۧ0��-:��F�qDH�ڬ���  ���.�{�7w�%����ykaI�j�mmۙ��H����uHv�������<�#�	B�U�����r��!��4��W5���v#�#<"aJ���z��`���h�l9��.��	��8������\K���i��4���`��e����t��t�S1��%�޹+|v�M�9�D�~RX<
)A_^�P�>=Q�#/qy>����v]�4�9��������Fr@IW@�hn�G"��o�n�*??��/�$�$t�k��(��fN^�C#����l�x�j�i�p����`ba��x�ψ˜V�gdh�+l�bЉ�V7�M�?�$��b�+���������3��Buc o��iuA�b\⸓��Y3c)���FA�rid��U �p(P� ��q��{O"�Z0�#�`����G1��<�O�1�v?L��f�kn^�lx���n��&Wm��7�vHEO���#c�t����e��l��l��c:�1����˶��"i��l��n�y)y2��1Q��I%�s��1C�L����~��Š?U$줠����(�qJ�V����X$�n�A(�Ǜ�������9��V	�!���k��vy���s�x
Ԉ��Qi���eF���
GX�X�F�� �
d���x?xvw}�_��>��~�S�O)�v@�K�:�O*��mT�9�f��欕�qI�W�����D��og�V�?ab��?�H��wIS��k&ۆ
d���b��1����b$����hy��X��D��?N���y~�x�(�S�x�.�ӗ����ۢ�)�w�����.M
ɫ^ ��8QA�Ы�$)��z�N��A���i��������
}?ߣ�O�y���:U-)����E�P��!^��rzwB�S�:V�?�%����ƕV��jJ�H��i��BZrs7�s�?�Z����1MlA��|�7?U�8Q)���+�<ݒo�j*K`�p8`T.gP+��#��:bݥC�G�R�(H�.3����'@c�s09�lH5�!��Ã-Ccq��Ӆ|l�%d��f�A��A)�?a��`� ���=zǔmٱB�1}D>�B�F��xF�s�N�pK���S?<=�r�_��t�Z/��}^O�^�n&^ _���cd��S�Tkk���V���P,z��@c_�"5�&�DO	���w���<�tpV�t�蠀(P:m��	bE��@'���KZk�H�Rs$�8��Tn�A�܈#����agW}�X���C��9��'޴��R02V:m\�:,��i4Zi������^/����L�J�G�3�o��7^<	;�Qs'NE�7\]MM�Is�RI&~_�J �Â�����s,����B��k@7���^N�y=̰��f]��I{+n�m9kY6���v0�nW$8���KL�}�XowwTc��e�E�p"�=L�}�no�B��OldǬ��q�\����ˉ6�eث�̚\�Y��Ê�qd[6̨"Ю0
�hg���?qP�'��p����6�	�v5�6�v�f�)34���M[\S�򀨿iK�\Jg4U�2	�yl$���UU�v�� ��pt�<1y�¨����{��V*�� ���u�M�P�A�+NĤH����t����.�uX&l�B�k_� |�q�+
�gz�q}ޛraaa�4��Q)u�w��
kKJ߁Qo��i�s$bp�� ����]Gp�7�AJz�1vt��ᎁ�"�y����v����0���hС��O ;M��.��r"UO����D�l�G�� �%HCeE�ȅ�/?�����{�B��v�6�E�ס�\_���	x���m�.VX�u��bt
a�d���E�౲)��~7%�����ѥ�:NDN�Fm\�~\d�X��`
���H�V��+�c��傒5C�F�>����ʠ�x�f�k��|X�m�ddc�Cb�w2��S���ԏǆie���h��{tJ��3�ז�trlLZc����'.�������wiQ~�YڌY�����]���JP�`P%��~����K<0���ͧ�}�>�&�;��t��Vr�|ij�%��g�W����H9��2O�m�7�'
m����DqO~N�n*#:��Z��a�e���]�>�;�_��
��@��*CpzFb�;��:;��5`�{脷Xh�g�� �VE�k�F�N"�B�-P��QRX���]V
��l�p�p�ɛ�8�S�5�d˥Io*��e�>|<e�^G�4%n�&u��,V��iqu�/��������U>~�?��\����sfW7,�8��(W�����Px�EFNd�ñ�''\4+&�
���^!/H���;�����_4R��q]����o�-Tr%1.�𬡹Q���-S�����$LGb7����aE��p��P��P���D��6�i�:&އze��pˮͦUJ@Gkt�\?e���`�}߃�x���P��Dt��P��a
@��\5��"��*h��:o1\[P��lj~WL�z� ������<�'~�J3ɚ[[���8���c���åzSP�]Q��ܽ����IL��t*���~�bU�d���!퀖�:q�ȏ�mc������"���,�T��t��;�道��Y�l��p�I��׼~�w����wg���#�6�ѭ]�g"3��f��K��w�S���gFР[���Y��}�PJ��o׼�~�ww�����H������<���Ӡ���f�{��G��]g9�%�f����hĶV^�p9�J븸�āE�I��5��d�2����M8Ʀ�/\2�f%�+�nV&83&���������Q�o��ǥSZ�@�O�g\SS
�E�WY(�.��I�Zݬ���R�q���K�=A#����5��)��´_�;�6�6�Q�{贮�q�/8	��Ob̓X�7а��nTb�n��S8$d� K�D�lׁC#mO���Lؙ���ӻ���Y��6]%2��TA��CQ�Oȏ��q^�ț�H,�6M��7n�&*�f�Aab�()A͂�������i^��S�����`Ċ{�������ز��\$��p��yzzڎ���{m�7��&ʥM �T$(L:ߖ���i���Ȍ=�����0T�ޘoI��{�,G���:./��Xr�}c�N�3 ���Ì[���R�Զa-f�*Ж����	��{wP3�����{l3�m�2���6��jg�n@hz����-�<e����=��Q�����`�!B��������ǎ�j�L�l�|5zn%�8&ْf��9vN�A������ʱ��W������YƁ� ���!S�
�ʮ��oƫ�{t� �so��k���r��:c�v h$V��Of��̬,f��+��[@�U�f2�+3�I ���(�4 -(�gP�JA��UWR&DF��XB�>o�рu�l]B��\�K��A��ʊ��|D-�+��l'�����E��]P��9|:r>=R�('�H`5t~q�T+6:���d��~o0��f��G~,��X�cH�������T ^!���,�?����Ǉz�����i1b#��p����M	�ۈ��O�CX���Wc;4�XWTx���XM/��B�� ��Ů����&�6�d�L���[z���R��TEF���kE����C��r�V�s{�K�q���w�SZ�	�$@�o���g���[D��nX���\��ܵy��p��h0��,lH��x�ĩ\�����]�� kTm����޽��]�Yo�ۺ33Shp�{��rSH����ߤ�1��,F�_��<,�Ne<m!���f���ώ `m?������n�!hK�c%�E/���O���=1��7f�_Z�o�+Ru?��*_ۂx�Դ�/2؎���\/Z��� ��6q�Fήj�t˗��|��w�hL%_)Pli�����-���`��و3���t�f��Y����Vd���`�,{������o#��n�3|ig�GO�Ǆ��oG�A{,���>�\.�&�ޘ��a:��	���w��ѽne�(��|u��n�"���%�n�c�[��aW���4a젶�:j���&��G��l�����t���I)��ʂ�E:C�X}l_YX�K��py�����ݜ�u?+�5��||>�Jml��2lЀ�o+��c����2:C���M�#�X�`���Ll�߾�7tN����� i�&Ce��iϸ�a��<�l�&�:����}M��|��h�si�U�Q?��{���=g��J>�r)!�a��=�K�`ac;����һ������e8�r��z�>'/PЁ�a�7=��4�3P����'///�ܥ� �j���zG�B���g$�}S=��u���9JM}����7�j@�-++��˝Ǘ���$H�_s����;=D>�#�kk�1S##%�or��P��;]A�2����?��v�$0 ����L�4.^x�^�s �B�
k�h��4sՙ�V��� �:������0e���vy�����m��%��k�K8d�X4���0���v�m�*1m('`7���x��|���ޱ@����XE�l���N�2}��C�i�	��P
ح��yw���PP�u;��&=��ק�]k ���3擤�����,��>A�
�]�벾���<�>�g���~�y����oȶ�>5��*�4��Z��3����8k6Z����ۏ���-Y
ԕ�wو�fg(�1�T��p֡3Э���Y8���XkӶic�3��DG�3���#�oƦ�/L8�w7��Jxo%��tY}�4ra�O<�FՓ���ݫI��L�E�VU(�_�s�o�O��q���d
��ۃ1����Lu�� Hx�@�� t9=W�a�ˣ_e��d���RC�qf����Al�;P�gf��`��PȄ�ې��Ǒ��-��S��w\ȾO�rŎ��v���ώOې�:�A#�i����uG�
�5^�-�Pcxq(���^�T���%`��zSj%�k=�&@W��;V���2V�d�8�u���g>������c�?ܛ�N2>Kw�f_} #2$$k�3�"���e���y'�b\� D�7*F�����$�4��v6\�.�P�BM�����Ƚwéj�utu�.����s�4�����#�~@������d2�5������ͺe5���+V=$��1�~u<żZ��)����HU-��4�4�Q�i������vFj�@ �/����V�Ӳal�f�6���G�~��ir]��O|,�4yw��P+����]�ܾD�p���u+ٶ-�����ԏq�њ����T� �n�&S���^;����G�2��`O���#W�_�<:[+�(�N�}C\�uۅw�Z�˹�H�h)��m�)<�vm�2�=�3��Λ�?��IQ�V���阘�.h�3o흝���6�4��v���R�mml�q��c��VVh�gwI���5NP3Q໣�RF��W�J�vYGoX�4���D��5��҂*L�ۆn�v'�Z�Cl��k���V�<k3��}�W1幆�ڏ�LLD��j׬k]��x�ƚN��C
~�сEtw����ڭr���Wv��:�݈�9����'OML�"��_�P���^��b���b��^\�Ubd_���}���8���W�э��c��%��|�i|��z�4��Y�X$�j���0�ŷ�v�vEx3����03c߬>]��֤3 ��A�F��ˬ�{��ZMB#FI[b�Ա�^�Ib��<ms&��ң�x���G��nյna��L��u������� ��<a�Q8,��PX�����}Z�շ�M��k�"�sף�����S��i�=�����!Կ<�G������Rn(�4�$̩�m�@�������IDN݁yCAq��x��\[~�H
��Kv�����#�g#���S��Faq����^�������1�Z��<h+N�Gk.�4�>����!��՝w�|�\m3���(b�Y9GA1�8�6.V Z�6d��\���=;���!`Y[q����b�Bz��b�V!e�_Q�'8D7�����������N�l��m�?�I���j6�lI�
ǋ3fq���p�p1��v+� RZ��G������Bm���Fd�g�ӳ��_Q�RM���l�|��i���v�}���B�LR��
f��X��+�kRcR�x|���T2i�g�d������stGS9_z�X����Z�����R� 6���U�����R:`u(�L���
$#���.'?���VOA�Km b��~oF���Z���� �'��~MvQ��|�%����a�@k�Q�<�1'ڑ�B�49�D(��0Ӧ�mϜ��)7ЅV?]��[�i�@T�/5m�۽X��������v+�|�l0K�~.�{39?�p���O��:��瀑��9�?gF.�l�+[�MȊ�&�?q쮒F�Պ3ٗs���qoseL�gff�����i�#G�=+�(�W��:8u�����
��ȳ�Vl���>ÐN:!��GK;z�I�|5?�-�7�H��E��L�0j�[��tvZ57��
�0��^X��m�(3�;�n�����y����l�gSk��wgV���z8��w�b䴺�g��Z��ۼr���xY�w�h����+&�p�!ָlX����q�����g0ϊ��]{_�%��ު�|y,G��Cg�}�a�������0Kz�RƊER�3�!M��KY�$��T�9K~/C��`���ݲ����1��9�ud�1@z̔�����ڰ8IЂ�$�eb(��H��b�h�)�Ğ�̪7⌠�À�>�Z��(rޜ|�t,��C���R%T�Vk0P&�Xqal祅fq�m���/,��m	�)d����Fg)�({*��T	�y-��]��ea���>#���0k�(a2�}��2ܗ�1��W$P,))I�ً.9�Q�A�5d�>�6�C#�D����R����x���c���"O�������}_)�Ok��o��3���	@~�t�r���r�b�+�����H(\�4�АUI7�a�tβg�[3���#h]��o���8��+�J�|��xg6~\���#����A�b��o�ڞ`aɆe�%��֐��-��۝�聫��;X�\�y�J��U�*߇���B����ͧ1&9)T�V�h��^O ��Q���2"�SKYK�=��z8�n&B4�d���݈y�?�_܏��F�.{�rg����� B��i�X�}�$;ܫ�ό����ٶ�C2��u�,�)���F��Z�����S�P��_���;�������
���/�?KئE�?9'����D�M��&r��I�혍=jӦip������?~��h�^0T`���'	�	�Ť1
@0�^*�6$_n�޿:�)����Rk�^�z�O�AU�O$"b��.��h"����2k#���z#uw��}Dx^�ZH${�8�?Z,w�ʺ��fI�>��Vg��e�C;.V��`Q�>�l��ޠ�I����v�B�#e�/cY�q�[P���l����X�k�����`�F�X-GabO�����Z���JIV���[��pJ��(�3tb�\4��mNT44��UNl,��@v�젳��^�s��%���@���f�����m�唱��$H.��x$S��-�ӆ���������w��1�; >s��e���ri���z����Nd�ئy�$�i}[э���:�_����X����?<��ed���X;G�����}�pc �=��n
�F�"O�H�q/��>��%�/�:�ߺ��M)5]�8�l�����r������#���� �#p(�܄Z�t��4j4XG����㱅23�������V~G���i�5k9{�X�\ƥ8�3/��JZ�ç��_[ �7��'o����t}n"0f̓����noˉ������֕���K#�J�˷�9Ò�}���ӭJ���0ѽ�ũ��M�j�@��dߣb?�;y�y^ÄGǋȉE*��=;��{5��II��pEJEJT�<��ٜqUp��T�pt�o����މOK���}�[Sݳ�R�����Ԡ�PE�(E:�4)	�W)�	���ނ�H����B����˛<��=�{�����C>�u�����{���D+��ǧ�J�PCl�����١ZYݢ�Q̅���}����a����(f�t����9f�T�aҌ����&�s/�ܭңg���ݠ�r����|NE����g���s����!�;@ǯd4��o
��E��r�baT]֧ԑjR9@"���b
+��j[����{�(e4!�x��1{sብ���,��Zen�/{��x����KI*��d������77K䬢\( /s���S��(�#�b <U��0�0����<��z������8�W�uc�9H�RRho#����Y/%���y9c%,1F���c�[	��T�S
��=��� 5��)Q��]�V����u}??����t���C[<�[J�"��P����P�8²z�1�|���&h��3�-��fix�c��� �c��C%�&����P����UEQ�I�+۹V�\���j�v&/D�b�c��&����H΄��������ݏY[[N���<�bM�)1��o�}/��]F��Y� ���%Ě��A�K�<a ����9�Fl�θ�VW���Mג��$c��?Qj(0���0�β3�{窃 H� 8J̃��Չ��R&:<ݞ�hh���N�$��ց�kE�'ZY�\M���.ɭ]�i��,� �� %�k@ϒ%����rv�C�`k���2K��:d��2a�a[�F}����::Z��T5	d]���^ww����XSM���.|�r��1Zi,�m���sdb���O懆�����Kum�E[ZZ4'l)s�]������2�O��圆;��#�����Qӌ���� �[q��wi������)6����E�h�hAa���$�+�@V5r����)�5ｘ�As�Ǐ~$��,L��LI�_ʺ�O�]9�ĕ0����Ͳw=2l���n����'����ؖpD�����ߡ6�Z)�=�v��eFp�s	�eZ� �<o�'�;?]�r��)*ѽ����]�:���v2��(a�ǳ]՘�6K�m��(2G���ۈ�I��O�p ��JX^����\��]|��ݲ�"�75p�~~�@�QK?j�O�����c�CHHA�aN�t�������2sޭŃ�GQï�DK�5 :M�~�]X�o';�uo�hr1��&qq����#�j��Q��	�|���C0M2~��GV���A�nމ�v��N).����,5�-|J�%�TK�.n�y�#��_��-y&0��3�F�a]�U���{	Q��lS�HW��jnO��4>�@� <�"�\B(X�g����~�$�G6%�&!6V�"ge&M8�G����	�m�Ԓh(�<o�VI[���W+�=�d=��ܯ�ӄV���.��[�n�\_�''n5��E:𩙙C&K�}uW��^����0�Zҫ�9s%�L���H�����n���ƃ"�*ѮP4*;��`5��JP���
R��%#S��H�r;�Mv ��-e_l^5����V�"���9��%�j��鑓� -,,����{`���N�6|�}����[c�r�`�H"֕��vxX=���s=>��,E%�1��C�(�!,��ܘ@��D���y��J�E����Q��߰W����ճ����"�,_v���m�TC_���O�gމ90��8���w�n2z:��r�<fpK6=���>N^qt�245B���RT����}��NpU\[Ԏݓ���KmYci=���/{��{ee=8�S\���ya;��8�f@�&'���~�[{%0�8�����I9��W��I+���|���n�<���/�.:���-zB�7Q����)�D�$r��䞽�����p�x��k�����C�����6���tu������`>�R�/�KF�"{�� ��5��N��A�C���!!m恬�b�i*O��L�&�S����ow/��1�^vy���kY �{6T��P���ĵVp-?+:s@�dl5��c�X��(}�w8�#����a���P}1W-n�N��HK��W嫾�A %¬�:d��|�M�E>Y�G*�{�wO�iJ���s6���*�0 ��XZ#����]l� ��r��o��P�щ�k�׌��it������hN��?d�;M����Z����)gb����̖s�k�����mm���u�e���jSR��;���ߐ\���tH����Ϫadd������磥��w�?���U_���8�t{�X�+uyӬ���
�0�
	�� ��qp����U�*L$ũ�YX�K�2vԍ:w��[[g��$��!kW��0`ʽ�'1s�Y�`���.[A�5d���ʞ���/���QC]�Gt�۫_R��^��(� ��s8���!��0��TK�1���P�<0,\'���6�^�=:���F�K|�մm��9��3kn7����Ħ�X@l�xgj|��zH�YW�i��?(O�j&E����f%��},y^���;����R����r��T�V^V.�E��qw�p�l[Ʀ�
�uc�'�@��&�|j���Ŧ�'��v��Q�Ey*��~S��A����zXV��>���g�#�6J�rG�/��E�����=�@�C:N��t|��K_������t���l=��a0U�� )���:Hc��N������݄� .��lEұa尹���	=M�q��Jc%����8c�i�S)�m}T���b��T��`Lr��gP@i��5�q��$r��H�'Æ�� 8�%:/�66��a����8�7e�t�	[�#>�Ut��᙮����s�����HQ�s�##@�d_�tG�f��E��c^Ѳ����-g^Dw���9E�-杩>��/��~���s ǁ�U��v�C��?.�R���c�\or�p�@U���ɱ�
�`��)^��n!�~��I�t��²��j��YOO�����:,WN�#Q��k�i���V�.�`B���S�ﵤ4��B�I����?����w|h?��Ԉ��^�
'%p�Muf�ڋ��z�z��7n	6��S�?�=�n�f��<~��I��shi�>ӓ3SO�3J�+D�tZ���k��*�0���D���hǘ���P������98������M�mM(1{��U�	�0���v�w����8Ϗ�_����լ����B��z�'����/�+eMC��l�jǅ�/u�����g�g͖�ʀ�v�!��͛o�==���cC%�1*\6p��	j���}igYˮ|������0����T���h��_\�$	��
?�Y���� �/��A�K-f�K��/8��*��OIU#
���-޻��0�����-s��*�� ^P_���� �E�B��;�,�_	�|��z������A��* ���z�I62���L꾔'Ŀ��x.���vd��Ɂxttt����ls���I�y6�L�]Z6�"+{���u����:&��(�[H/�x�B�h�+Kk�Y�����`.�/Ù
������9�j�.Ώ6�Gߡ6��?ۼxM{1+��&`1~���K�����@h��[�Z6�'+��-Ǩ!�T��?�yUh�j�Wme���e>����Vs��OPi��v*��3��2�_�u�&�vy�}�lZbmĢ'��{�1HqV��Z?I�Ą�zσ��_Q�S���<�Ǝ���� ir\���o���_��ʐ�
@�QR12g*�40-݀o5л�'�~W�j�傒*��V�4d������2��"�d&�t�'&%m��|��{5�i[5|^�i�~ NBV�ΜW�����c]��׵�|��w�>�j����R<��kv��!͸��v�*]��9%����6˼��x6�>��W���qsq3���+tyD��˾q�		j2I��'��y�~�<Z������i7`��2��e;���q��*��?�2����hb���sѴ8MX1��|�=ok���!�$_����uG�b_������,��,:O�4�-o�d�����fh�z�����}vT�Rx�l�&_���Molp�ngww�~[�����(�c�3|��1`�4�d0�1g����橰�D��3&�P"6t��~���i�ȧI���� �ؔ�YL\�e����D�fhO�-���wL�d�^��0����2�F�=
}mm��/�	am�:����e1D7��kM�*F3*~�v;�&�p�=9>��H�"�s�)W�����@D��*�{�Q���j���)
�(�8��O�ea��) kPi��jk���J�4e�M�PQ&i$�B+Q���tGhid2�yҬ*�b|b�s<+��X��!��݈���5Ɇ~gdۣ�P���Y#;�8Si�*�� �w+%/�ɟ����۠,�#�8�F(\���ӿ�[�f�Q�׽L��o���嬗��%oDu��A����o�9�ZP{s>�`#���˶B� �,���Ϩv���\I�p������e���2|0a�܈L�3!?�"�̭�:�<��i��b���C��zS�xѺI�4��Vh�֝Ւ�qQ�jT�'����_�>+9��J	m}X��B��úYcV���brCC	�����2�M��~����GZ�3�#8���m�SfP"� "��-iv�7r�Zr����������en�$� <��{�0�n�B�n�Q�M0�������M�B�"?-���-8�Ս(SE��H���b�E`���U*���x�)�7��x���y�������Z������ʒ3�K��=��V�<����S�P._Ŗ84���e�Z�(�8�D���&�gҘZ�B��������1u�����c��ҐRL%ך	�����'b��no�nm��ģk��o޴�Mo�SI.�6n���iaq1G|[���[^�E����k��ʫ�+����JɁ�-��s�@�)9��w�ˎ7�E$R�W��ZL�iB>1����|���=�1��oﺟ�_��4#-���O����xo��P}����1��''�v.�/_�������,E(^�V.���ڡؼP��*�p1Q���x�j�ɿ�:)C�����`_/5�FK%ؾ/^�jL��ɡ�S_�>������M:��^"�3ss-�K�.$���%zŗ��}]ޗ�1P�YG`��@,�Yz��+���ܣ�������+�}!���F�_x�&�f��*�i-}�&�s�1G�hT[��yy��o�Kf1�qtj���d�Ӧyu�C���y�f,u]��i���g�'�H�:n҅�)���׭R��R��������?Px1yj��*�5a���$�9����%�N�8��e�덙�RL��1}��ɳJ�Mҟ���$RY��sksg��������#O4�'<���{���t���%��M|����J�&�^ ,~���(�xQ��ht��E���zR�l�C O�JJ:�h�<C�Δz>��to���S{��.�`ݓvW7�f�Z�x�}����?k�굺�70p^�!��u]Mr���/d^�-ȳܘ��q���,��� ӛx��RXXؼJ�+)�]oe�ZӞP�C�1O�{Ͻ��z�p�,x�Ĺ��WQi�*uյ������	�+Wċt����%��Ml�g�to�ٴzp{���p��'��2/{����4ߺH�I�\�#�p���\�r#`&4y���ˁӤՒ%�Y�ʓ�"L�a?%[�d��"�2�Wi�n(gd#��L|D�O���_��;Td����� �%o8�oo�W�r�YT{��C�-s��Y�84�A0��J�zkd��"���;W���P9c>��Ծ�����M,�^��PJ6Ϻ�u��_�HH\t�@�sKdqv�$�r\@81���� T���=�kW,a���˛�p�w� ��,�������<Bɳ#����⟦+�I��G�` ڽ�D��L�[�c�r�I��v���e 46�1Z���/��VDT�U�rn��`蔡��P,H��=1�y����C�����y[r�b���C\���W1�=>�خ�t���ߞsxl����-�U\������lq�0��U4/*]v���,K����U$���`�U�cG��Y1/2qŢR��|��[�'p����g+��t֬��b�s�.��I���$.K�B�j�W|�;.��;������tQU��9�fE�:�J��AG^���pq*Q��<,k3�g��D+�f�� x��)�bP^��Y��H:�7�@�\4q�qy^Om���$O�Q���m�X����\ ǅw���w�F>�'��`<���S���z�?�"��\&��'��(���T%����)�^��Y�
صy@Q�G�(�/��R��p���J�4�6e������K	�]#�-�]���=n�Jyd1;u�5�=]��ovh�c)���\{K����ɳ�3�' ף�x8p��A,R>���R4�boo_�Zb��c��&������3�>�Ж�L�x�q�=~R�v\)���Ȱ�3XK�?�=�:���{��D���Qfw���� Pc�wA�M'A�5��ș�D�X41�Y����?�\P
�}��"6��H���B��b��m�:�ox�	Vb�����;�Ǖ�@���J�����׭�p�U �%�8	�MC�?Cc�tƑ1�J�%�8	��?C�6Xи������q�D8�H�&�5I\ �<�������jl~��I<
Lé]2K���*��?)h��6X�'Ѥ���[؟����ϗ>�PK   �	.X�:sJ� j /   images/920576d2-9ce5-4348-9cff-973310077ed8.png4zct&M�nrǶm��۶͉5�mLlNlsbۚ�N�<��Ώ^��k׮��VW���$,.,����
�Կc�ߝ�τ�'PWIQ��i�3biq5O��n�}�4���FLm	�h����b�(T
�ݢ��B!��<c�<K���^;��z��A�Rˎ%����h�9C9���&GN��#�;��,�ݒ����[>W<;����:>�%��2tJ:A���~�.�4J0�k��!�^1�A�����B��FW�xB�j���˞�_�V@	��y����m}�M ���؞���4�_M CG���媇��)��:A���@C�3%���O��}����_F'���;1u���/ߊ�x��G���Fo���QZ���y�������m�T�O�6@��r���K���v�5��@nkMpv�����q�^���bZ��<�p���*_&�ʅgN�i%���ϕ@�!�=;./��])z ��;�S�����ߋh��4`@����5<�������f�U�����w(�ϟV?��mO�Q_��Ϝ9��`��[�'�]�{�通�`�K*J򯍬�ܻ��#~�0s樂6��r��Ǻ��'�g!J1���D�(�C�k����f��f�Y�т;A����q�\s��1[��5O��};�<Fb\m���eR|2�uQ���ʭ���3�qT�_�H[�P���m��"�e�t��U�^kO
-��C~��}�A�yp�^l�'q���Q��X�;�s^��Ps�;-S�}�d���	
l����[�zVY��Bus���J6~�+۬�X�I��JF�i�������D�-�ğ�ƿYj���j~��4�;<�e]è�_4>;w=H�|i�y��y���Dy�~�2��S�:�����X���
�Ќ��¬R	7���ڣDx}ɡٽv/+�_�����'����8�r�}3� P)}6�_C�_�w?�g~��r�uT���g��l�X�Y��J�ۃٜ�9Uܳ⏊���:��f�\����AL4TXa&1l����Ǌ٫��<�k�η��˕W]�O�8���{�v�y�oi�}�|%tz|}Բ������d�'ĭ��ʲ���e�%��S���XȔ=�v`.blj���~�#d�����,�[�ctP��jU1_ 	='�RiS���G^�᥷n�{h��	�'`�h7n�X=�q���Z{t�?�%wm#(��kl�����;�G��}c9(d��mO3<�NKA��)��s̱פ��('%�1��}��ԕ%�Z�,6��y^m�*��wՀ����o���]@g�7���i�_�<�f�M��^��+Q�߫�Y9���N�2+�T���/=@7����[��,��ݱ��Mv"h7+o��HPɅY�U����Dj�����L'}�@�a��'�`��E�Ch�>؈%�Y�U�7z���;J<E"5���)��H-�N;��D�py�H'"`%y���H�r em�U�(e63꘦��[�h'(d���v��=%_䚶����e�汫���M���+��	�W�X���^�8�~?^A͓����T�L���,��d�_�R[�|$"��-P���CDeA��*AG �bf� d� ���a���D|P�*צ���J`c���F�YCծ8-,�X+2g��z��nۮc�N��Q�`~�����Ka�id����~cw ��:ka2�ϙ���"��-Nn�MXq�z�)*؛�.��W<�:��ƒ�G��{?�>���˥��m������Ĺ�۠�77o���՗���[>����RJ�=��μ�'���W�"Q@� �$� ������/�"
8.P\�t)F�V_�ڒ`�A�x�Vk%q�u8�9�O[�F-�F+�>Z�^�`�W^�;^�̗�6�� ��@�ߑQ�g�^)�K<~��A�g�S������3�iÂA�p�8�6���CVT�
�����;�U�m�{qC��w���i�.�w�B�|������R ����Y�������[d��eEE"g��
��+.�a2;�P�Q3�^ie_�:r,��y�V��x*����,��Փ����-W�c>T;��9Sb�53�a�W]��!�i<�@���P��C�Ș�g�HHs=���/�:E����b|gP.!�D#��؀*_�^7���
W��nyw0)[�}c�
е��P��Q�bɦɧ��#QU�tT��}N�\�/����s�!�����Z���ct���ѺO�
r����3CT}�1�6��:���G�{� �a��/�2H7���F�4_~+Xb�K_X-:�@E�k#�z�r)n�O��##�u�)C�V��3/�:�L���v���X?}�dP[6����B����|���(]��jgb�O<K>��+>�Qy%�<O���B"���V4RJ'�v�HP/$7�+�C�Y,�P�J��_*��7P�l�K��zzmv�������VwuX�U���nt=g��-���[m-��6u� ��'�^����#� ���!"����uu2��u�;^C`�+�#%)�J����$� �o�`�̂�0���m����h� ��'<��&y	#�B86c���1<�h�#����H�)�e2P������[�%)�Q�!z� [	�K[u����Ae�^7�r��`������ ����^���]��8��KVoae�7��nN,٢��Tm��������y�������2x�Pqb�5�4W����.y~�2i����}��I����=$�M�����<�K?��9�G�j`i,H�j=r]��z< Vj�2�@���&%�O���O�iDl���s�("aF����;�����d����5v�.��1�k�hŝ������⢻W�g�U��Z��X����������cJ)�V�D�+��2(�I����d��Qآ�M��ee�'7"(�h+����FÆO9o��ƥ6~�B�ߖ���%����.��#�s����q����Z��ٳ��+��N�OЎLT����c�71�շ�\�]�o:�ϱ}����B���Tb�"������v����*ɪ�|��DV���,�{�#�"���.�!��䐩YC�%~-����5��B#�@3WF2��R0y�,X���솹ɻwhU �W�kB?���r��\���xĘ���|���I�S�$�Ü'���+�
�A�-��N�ˁ5	"sVn��5V��������"~Diƕ˹�%󾽋�㳮D��@��-�n�@�4���DF�e���sꧼ�K�o��4:�P	J�G�ԥ��ʿ�;�V9~��_Y_>W����%�D��) w�/��N�����g���y'e���*hy������?���)����� �l���bF���(�}j�}�M�s���I6x�*�w!f��	��mD��)2�R}M����D̑�உP4}U}Z%�5Y2�{O%s���<��?����d�� ���@��e!�G��\7�>�e�yap���K�H-������ҫ� %��5h�Ρ��h��UL4\E��Y���	����Q؟.�`;�����Ŏ�8�,[��m��~^V�z��=�����M��0��q}A>�z�6ygB����\�檭}��]d5�o�o�P�5O�4�֓:��@n�� R � x�ӘUQ9�T��*��ݒBQycÒ������r�Y�Sʮ@VQx�h`A6f�0ɵ0�4&I�~��!ZH�';�B�����ڊ���S�@L�Q_�T �\;Ѭ�~�G2��B�(���B�pr���D����	��@߸Ǉ�鋨� �^8t>��;���	:��<�V�Z��~�<@�Ш=����|�7�W�����Z��#��1���nK-�4^�7�������r;Q�v�SV���@|�o�GD���j�)��
��8?�VŔ�w�bcb�+����J�a�G��?W��\���7t�y��AY�|�af��h�"h��n�_��\�E +�����2YĲ4��oʰ 	(- N�6����}7�P`���疫r�#ǔ�JɐV$�����
��j�] 4�g��'$�H�t��q�T��J�ܒ���`D��� �X�j�"~�H]��� ����²�:n�q
�t�;�Т8�,I}K�;*5�7f��1a�Of�	!`/.�A��g[+~.55��8��cY�a���&K����k�ٳ����x��tN���U�yޢ�O�o�����N;�0[n�]���������*��+�[Z�Q��P[dc���N���O
�09Z�[�%�(�,�h���YE�L[�+m;Z��z[[}��c�,Y=��K���R`1�_�UC��R3�(�8kԛW��[_?)��5c�q������;r�`Y�'S��U��}�Z�Q?��N��^��T[� �6��⏔�	�����#a㈭�t..SU	���v7AҶF���ۉ�K̒)GJ�;"��"Z��i� U`���O4�U	��G��6S��ҵ,j�#�����=&�x0vq�_I��G��6"��#`dOҩVn|L�6{p���A�6���E��8G���=zڵ�4tzM_<�����k�e��<*�Z���8)4{�"xl��w�!v�'{�S��ʳ�K)��^�f�l������sn]MYK*��,f�^�X���~̠�Hg
�u�H�c��B6js��,΁�_�C���l�eF��?#���I�����+=J-�x�މbm���� k�X́�h4�[�N�?j��`����u�_L#�.�!'�Ah`j����WsD�3�{�`�s�;��O�{����p)E�Z��qF�EJ���̺��	l�vx�&]$��F�ЉF���|�j;ϋ]m;3�Um��5�	��R<�{����SO�?!cp�Pkϊ�[��c�n{�.1���<w�k!Y������킭ɘ��x=�4G��t�$<q�A�fܡ��;������SPA�L�l�"�:��in���0Zsy�c��P�]���^%�����&����w]�`{������3�K�������]�Oc�jS��d��Yq��U��(��
��YV���N+�&-Tm��>pzY)���Tt�T,>JJJp�Q*��E/��N,0}�yc4.wl��A�l#�Z���^sw.Vi�lJk�!K?��:�X~\�GFu�~�����7�'7��L^�$2�7�R���jb`�tӴ�`��}����^�}�o?JK�.yO�`6��6�[@�`����8�Kt&
�1�}v�n��hQ���Bȥ�Q�z��/���*���Jv��z˛a��WC9l9Σz��}���)V!���;����~����X���T��+���yU)̂�A�
������BN�ƙ�V7���]z.�hmG�4u��v����)�����u6`��������-M�~�e=.g�k�[�=\n�w:�	6K	��j��0��H�CS�w<X��:�E�O�=��1���J�F0=��tZM���Yӷ6b��y)���J����m�t5�EW�]y�%���gn��vn��u�ix�2rp�������5¢�t�ml�mE��|vIا��&���xf��,{�����6��d�Y#���Q[�%��c&���*M��㩌N���/�Z�P�l�Z��-�E�d��#���"E���
*Jꢂ�\�s������
��G3/3$S�p��1ߛ�:v�Ql6��6)��?��+���-�-�,U���#T覗o�����
���pX��!��E�$��� $�^���ω���Vj�z�GFA����|�
�[��M�Zǌ�軉� O��H�sί�j�{;��5�oȲ;��D��0��Q�n�����|3_���76S�@=.X*8p/lޢ��LRV7���y�4�*hS�ȶ�jjX@\j_��������m�ϰ[=�y��(��&��1'?MR����)ڱC�ǫ��X"�U($wWt酐#o�"6�����GV�'����f+�Fl��rGk�m����Df��\*$�<�W�%%��<��7A�r(
d�+�u�IcЪ��9n��D�4�Mp�EXi6dE������	
�`�-�B:��,4K�?�F���s8[�r���DO��	�u���}��V z�w�!��!@�R�(�8ƣdZ�':��c�Z���#&$G�	�!�?�8��������J\�
|'�@�,�
P?JƁ��4i�z-�Q�=S��5�Ҵک��y�����e!�R�_��+F{�據�VW�t�]4�P�%�����.�`����\x:��Ӈ���n����δD!�������6��q�@r���4�b�"�'9���	��@O���QC_P�e���#ٓHY�2��t��8���I������(�l��.�&� ���:��Ľec�FEӀF��k���e��; н#�n:Ȟ/b `GT�Dԏ'��Y�C�s�Q��|@AEme�t��r�͝�&;;HJ<���[�T��j����t��`^�fDD:64����⧢��L^�چ�]��N�=���N�(뉗�]����׷@baL�r�Ǔ�d��������aXT��=D���h���� ��+�
/Iz��=����^��ђ��Rٰ�܉��ӰY��*C�K��C���|M�ɨ�/w�u��R�h!5u��A�c!�J󺩒�6�å'�<a���r���Ɣ-�e�����l߼�MaW�<��g�g������ٓ�`Q4����{�À2��n���)��.Hٕ������I#<L�fDL���<���u�X�h.��J���:�Z�m&�,{x�/e/,=��H�Ѭt�.�Y�I#&I\��ßH���KUJ[Z�g��^�<4�IQ�]?U%�v5�>+@�U� ��D�G�VK�q����bV֎�'m�JW�YY�;�x��<�R	v�Q#i�!Teб5X˸�K"���\*�k⬈��ݛY�x�ۨT���1/FD���m0�oMG��,�;�g�!4��)�Q0>�fۄ�ʰ��].�b_����q2I�Y��xj2�ek8�!9���ߤ�$��e�d��a*t�)���������5҇�T6T���4�ãc���1�QY�����H-o�[x�k��<�[}�w�1�F�fs�����]�$V��Y�ՌB\��Hb&�$I~��)����� �9�Q��R�m��5��m�d��ƒ������+��fr�1�y��M��<ܠ�۪�^�*M#���()E���W�>�B�e��ʤ�ұ2֗ӕ����;#VB�aW�kv��z��&G�g_��n(�GФ�����d���l�أ =вx�~��7��kL�ơ��{S�?yl�-�ǵ|G�exI���RN�4�{�<��\����AS�WÕt�;�:"a�V���w0�Wk�(ܡ����;_���yX�j��W|��^��I:m��X�Zg�G�9�jt�)PQ��XR�]��ӻ�X�N��<1�;!%�������q��Ы�b�G��G ��{��r������T�Y5E%���}��7`x��Y�c�1R�D5�]��OƓ�O�����M.G�h;�����-���F��b�Ŷ�ds`��$/��^�!��x����}��@�T<⢑�����f8B�ô,d&Q82B�暆Hl	M*�^������n耉?<�	�;,.G�FQkۯ�&H�E�WbuK�ZK{==��ύ^��C��C��$��`���pl����M���Eh4��\Y^ߛ�u����ۢ�s	Q��6���®���)��A>�g�$�(3!'�Z8�l��౼V���M"��G*f�93;{���h�;'e��G��N�n�����+����?��0��i7��ަ6�-���2�jǥ�A;jH]��J��̴����5t�X�پ�?�� ����ׂ�Dl���;'/k`�������M�+�"e��Ӭ�S�ib��,���(�9�!��\ͬ\�3�=���_B��k���e16ZX\���4t�#�ɠ͙��wv�nh����K��s}L��O1�6�W�+��w��:=��}WZ�-�X��⁛K��5��C�+bS��~v'=\	j�q|F�0��~�)K�\aHU����l�Se�H���z�����iI�%h�譕���g��O��ũ	�@� P:1uW�G�;҆r���h�����������hF2�" �Ԇ^a�%r��呖��;��q�����8�H�m@	_� �Aظ`��������}v�1�0��fA
��|<��e�7QiÒ;�,.�3�.7���@��kgu>����e�ۙ���^�G�P~j��H�J�������5�v2	UD��S�^�<3!� ���j���yz�����h���v���f1�KUi�FN�R<��ϰ�yv�c�\|�A��+�b��.��2�+����E+	>sFI@ɍ(e"�]��N����SH<���>q{aD�
��C�J)]쩭���Pi�Á�g�_�"5:��}����|��x��{ĥsܥ;�\�O�����>��y���h�re��2����R(D.{Q��l���?��	��D[�G���.�<�-�IX�'�i�3"�$���{P��oI��#�.�_b��xĢ����� ftn�*z���5ϻ�k��;��y������|�\� �Q����3�.n�7Sw��o���!���[ݪV�Je�mH�XFV�d�.E��S�|��
��b\1�I���W��LKe��@tTټ�E5\K���������1�y!���-w*B�;��v�\OVW�RU��ޠ�d�[Q��et�F�� ��Q��rG,FQ~?��}�թ�W�N/H�h#�o�&1%�Ӻ����_2�7�g�����hh/��df��&e�u['8�9��R/tS�$��͌��r
Uh�h�؇����"�	y��{d[rzCOv hCD�OR�ms�|GV���9���Osm��嫬f�����g�Ë��~Z6��\����:��4E�0��N���[RL���y8b�)4mi�����b�/�"E����@	��0a�%��$3Up���͙��J�a7��'G�Bo ��z6���қ�K��D4�{��f�4���Ț,�$ň���6<���m�Jbk�h��o�����~Z��>��s��ďbΌn�׬��^]͛��`k���=��9vz^D�6ح��&aA��r���u�Nr9ݿ�W�H���U��V��-����.�I��q��������<���t�m,Ċr���61�J�ރ_��8�'c���	!^E���5�g��_���/?qʙ��̓:ϮlEww>�O�V�5�gs�\�1��L%Ȕ8/j_|�QM
!��K���0n���K炒X�ɕd�P8�
!�9�kO���4c(��U�D3���1�������p�۠�'qQ�9J�iU$�¸t~2�'�'�g�`Hg�("�,s�l5�|�ۍW<"���]����g=@;}4�N�cCO⮾�o��$)G�'���y^؍0��H���⦮"�n.���4�"qV��40�Y3Q�q�}��N����XS<x�(bF�Σ���'sM�`8�+�v�m�c�Y�ܨʉK�HA�]� w���y���
k|'�w�O|��ڹU�,S2�HR���D�hӽƣr;�����{ PRYC;T���|�QXB"��
�-�H �+�T�E	�8���R�|<j�����t�e^m�C̏�g��G�GB��k�S��8����ݦ7�-]"�j�>��� ������?3�%�n��"�B��b�'o#�Lb&��[J��x)�|qy9�X;vދ�\$pz�n�ׇ�����Ϗ�}���m�潔�)�b�V��سR ����<*�Y�o��t�^36�Z�'�Y�����]Tg8�Z^�	�؈�v�@������ +N�tcA�:�r��C�DW����u�G��w�����n��.q@|���5W.�����l�w!�v�4����~n9����9Ų����3�fV:��4�__��C�}�Հ�1�G��-�YH��r�i�A��+B�;�RH-�qC~����{���3y�,'����2����Ñ2#
�CsB8�.)-�B4y�D8�ܑ ��I��iJ�dy����K@S�$+��'k��l�!�(�z��-6f�V$�������
1�`h.Q@���7HT�/� C_%���v����d��1�
X	����m��>���U�c_�$��ύV8a=ݿ�]$�-L��%ls�r}Q�<f��'|M���=��F����$���HcAh����ʕ[�U�m�1�,�'�T2���8Ç��H���&�s�J�X�\(Q{ᲈ����"�m�C�� �e֎�%1u��P%���k7ZN�\3t�,�0i��TNU>��bP�SV�$V-ϱ�ھw��-��Ϝ3-�?��N�L�(����#Xu�D���SIq�@d�=���m+ i��:_A�Ye������lo��3�y[�p� �����U��u௰�quy4;0��)�c0a�c��5����ܰ���e\qΧ.i�K{^0��-�ilMќf���q���=�E�͔�6�P�[�5<�/�N\��N�T�ƘT%/1����r2�T�	\�G�$�d�v������Cfj�� z���j�h�r�:�B�%U��%�4C�3��[_ ck3d�h+�~�H|rS��I�I͖�xd4<&�����
�9�b-^Q�z�Q/�b���`��m�=�!�z��g ��r[g%�}�1!l�/5�QN�q��hyW�QL��79�)D#��y�����n�.�N���E9�D����%�����7�8�u)��dvV�C��}c���:,+�Z��5s�浆%�{z�q�;��bӭ�l#��;I�5tNԽ�Z5R�
V��m��k�:az1L/fx=�t�s|�vv,�f8\y_N�V�9<NԨO*���O�f�~������`׬Q{�2�u�L9�xr��L+5~��'�˵��L�D!G�����GW�a�����=	F
u-B>=|����aݶ������8ol��J�ŻNO9��4`S(�\5Z�f�Ο�^�,��8u*R0�%��#l��n�I�������@�9���|B`Қ6m���;Ʈ��z�2)o%r�ʾ�B!>�q]B"��p4�Za���f�I�&T�4v�z*Ȼ�4�6_����@'�%�L$�9��zO+9
z0���O	���֬gm@[I_��&��f��OEz+���Dt �^f����o���O��lZ����w�E��4��je̶�DOAe���ךT:�������'�{��T�1��FT�/���(AnϝdMƼ�:6S�tkN�2�ɛ�c6#n�	w�;I�9���+�m8sjr�N�&Կ{Q��ܝR2S�}���ñ@��Sy1�.�E�<�}���3����V9\����fQm�����R������W���>Qq<Fo���f����N��GFȃ��[�"M`<~���ߒ�Uɡ�O�z�6k6�\�4�Z��R����3&CWo�]�C₠�ݧѣ�uy�Zq���߭#��~��wBz;J�L��x�	�M�j�<~o��6�������I�8��b�w�v�ɺ]�#h�.��[\��o:'N���O�$��A�@���u�)I��?�VV�w�9�\_Vj�6��D�.:K�{���o��P��@�m�.����,����-Zg'��YK���R�.�<�0��f5EQ�O�H�L���
i�ӂנ���kGKeޯ6���;i�ksZ���ٮ\�oqP�8m}-O�= �n:�i�D$������\�o�뻱�B�XUӡ��C�G�Z���I9	9k��������4���Y���Y��CbM�p�"��m�X���"�t��j��!�L��|8�n�|p�/�Kf2P�K��M/�T4��u��t�������؜�q�Ⱥ��"	�uo@{���H@V)=��3���-��|�8|>�8�\���ޏT��'^�g�h�@2n���%�m�#�O,S��De��g���^�վ�p�\�G�:A��;�';���UL#$�1
�X��=_D�nDԖ��@�������}U�6u,9*F�F[�[�<�F\�ͬ���u�q1��P���({�k#,�M��s-g�g��O;<	8!vZ(tL;�c�1��x3�coO�m)m	����-�e��a�<a^���WW����5���'elȾ.a�����"a
��2��Ct4���vW���
�]DIG�s�*�̶ �k�:�����ȴ����P{A�z_�'�.�_�F��Zx2#���'��:�5�Y�TK�s�����=FBPJq���C-)$TĪ�i��gS�+m���䖳�?Ǉ��I)P�h�K�.�6T[����e�X�8u��dՔ�W(謂������O8�Ƒ��PVW�5��O��M>~�H�ΤK�$�P����`87M�ұ�(�<b��\�:)�?D�m��*�-��� ��������w�88o�������L�%7�^���ZҬ7��$FM�f�U~��=ܓ˗�X�|��P��fFB��Ź������;V�omc#ޏ��^w�Np�������
����p���9;L/O�Z�.�D�׿�x��C���Qg���n�"�w��>t�	i��xa5�ߠ�$�0	��ϯ�����gF�z�i1}~�'hK=�1C�x�O5���8D��������+�9[%�jdH����^K��5�]�|��6̘c��U��z���Ӑ`R�ckk��΀��5E��U�8~�f_\����Õ|m�\��X��3�E�0����;m�7��̒0u�;����}[�����:R�KS�TE��M�ES�v��K]�sҫ�Y�����@@�f��:��ͳ��/����u���k:_"��M��\Z���}*/�I f�*���E'V�MHbfȔ��m�37Ƣ\��0����0��7�И|�Ց���#�غPV�q;�p���
^���X��rFd�����*�oO�z�E�)��p��� ���~�cak�Eɰq5�v�d�wW���7mQ����L�q��n[<J��L��0�:���@��Q?"�_�5�^����]���!�S�cv����W�uL�'��"��k�Eo���z���5�a��)����D���w��B�0^~V�iQ�я-�L�"[�%u�dwU�"(:A�~T<�I�W~N���ڸ���J}�2���8lO}y%����u��������Qw!���MDv?J"�Ϲ�] �%V�^��I��dc9���Rs�a��g�.VW��P�3��SJ��Z$�C��0�3��p)��LUp��@'��Ss�u�|�����Gi�Sh��<w��Lɰ%�;�LZnv�?���u������%��= B��$�d7��}�_�e_�7�� Ă����|�mm��}�ɝ�ԭ:����*�-��������������^(�D�nнg3f� S�z��;^إ��iU��=�Ӄ�IYt���Pד�~�뽻�{�$E��e:_ ֞�P��B��<tHc���
���z�2�?�l��}���)1�%7,�,zP��t��X=�>��%�� /|;��9Pix���5�V�m�B��7������[�(��2�@Zb� ����QG�[��+؉�qk}qx���f ��c�/�|U��:��D�1��A��W�Mvy�߿F��km�����ͭK0�l>��縷ӓ/��"�V�`�{�����q�]�U-��r'k���5��Y��b�-�L(�L��@ -\y���=��"����<CY
��(m0<܃�4ź�5�Zi#>��i�/Uҁ�c�P��}��B�ak�%��J�~^��rD����y���+�0e�_��,̼Ŏ�Dǻڈ�!j#��dH�*�t�x��g�:��&��h��kA��t��s�:�
Y�$�XŊ���nu0���Bl�qͮ,��&S�~��m�dU�]	�������0s"
��ܫB�\_�ӹ���YXcc����WfP��,�
0�|+G��/3NF��� ��U���ң��:	�Ըr�����~i�ü$���B�Kj��֡�(+��W8sNW��lѓ ��V��.�?�hRrȪ�;B3c�c7J|���S���JxaR�˹CU�N���|�sρ fS��U�ڮ�@c��x_L�Y)��eG�$�])�P �ph,���' f��1�2��*��:��lm��N�w?�'ojK�K�x����?����e}xa4��%�F�Q(��V���o��)��n!,%��2b[)w����5��T�nf��=���ƕ���De�=��15�rܔ27x�!&��`��p[�s���f�Xd �*��B����E�����L�!�pv���\�ʀ�0�6�7��Hn]��������y��H�����zT^W��O����4��tlR��z�_Ug|���|�����/��+��)�-��<���b������qȕ�;�ӫ���M�R)..n���?�mTQ� iWE� �����k�ʗ���(<�mo���͎*�����@n�����+�qS�D�y�	��y/��
�jr�@���sa�yK�㑳&Ť��t>O��h���0\�*MŊ5v�ܝ�TI�	�iTU`1Mt�yT V��&r����.- ;���m��G�'��5EI����N�v�!�]��h/���L�*Rٵt���i���<�<�R��U�6ӳ�ov��;0�V��}�F�Ğ�d�8�7$0�"���&��p�EdU]&�"�d��\�"�%>�_ţ���*�*��NQ�
@x9]l�,����;��h1���\Tҥ_�F2��e�c��8��Ԋ,%�7�ÈO&k�S!���u�0w�aB�!3�]�ҥ��Y�F���`#44�T����1lBր�YI��/{��2,�-�S�e�!?M�&ya�KP�r��M���t:@k/���|�i:�v�-T�4{���`�}���e��P[\��Υ�O-E��q��w��-�����@���&2-���%w����㔥A��啕���J;,��a�@Q0���X&*�v�`�\�lQ!��d�5m�:&6��C�p����F�ǌFGW���7,�i��>w�YHΉ��7#[>�:�~�#����.��I��Ug���SA�1*ﰊ��R�RsP�8c�0;g����7�W�Z���;k"���Ϸ�	N�/ia"st��G��%k��*|����ms���u���Lj�	��=����O��w��ߒ����!�cދz�d`$�V>�����ĐTM�c�'�T��_��!�`�ۤ��t2�j�*ѹ:7t2)@���!5�7cJ�<�MW��9�f��@��>\���t��8��33+�դ���V����e���	��E��#�-�t=�Tڌy��d>Ҏ��/��*�ڐ��\��V�P�R��&{
��#��ߵ(;ʨ/E������%��=�>`�����7"=��5K��i8}v�$��$w&2.���W!�;h�*~��k�ý�;��j�eI5W�������r������42+�����Vr��B{8�>�Y�2<4�>22r��]�Nɗ���v4/1����N��Ř��S������P��+�.ΫZZ��QI�m3��G ��������QN�CC��'��,��_��N 1�PI�u��"��!�<f1^rN(Ŀ���'k�K��O��T��+V/w��	�	��A�Ś��;=����*�Y��ح�}İ�� ��W;Y!�y�3,���*-K���d}�=,q�D!$�����T됄uۂ��[L�Vf���)XU1�� �ʍyއ���D�B7�*��$���ɾz90�,͗���Ǜ-�zz��ɒ�S	[@Ϫ��k�l�KU�������P)k�e�A�ON�<2��m0zw����m�́A��w�B���3��I�V���Vh�$��ޱʕ������_��&h�1q|R�%H�K3�e.3%$�������M��_&��^����[X�8�2Ys�M4�?4b#�1��;j�/�#J��?_��'UD��\T���%ge����'��1��Y�?hd�dck�,�J���ה0���O.�f_��v���L����y^ۤ���Udb뫂y�+�"V����c2�<���<�� �{��-�DN0��[o�I��� �|:F�ʓ��z_%���-z�Z{_=����_r�y�tي���A��f�����j�����oo�qs"��&�����)w��i���|�8�e+�M�E*c]��L*�U�ut{�s��:�+��4'���J�V�hkIK��G��5'�꥟5���y��� $�� �9@�V���wF\��7Ż�uؼ�T��*�_�2���v�u�)�I�%ks���)$�~���2@Ϳ҉m<Y.��g���g�2O���©38��t�=�/� �ͺ�D��D=5��Q�![^x�eq�IB*��S�=���7���А��VT�$@D�	U��2�끇B}�,��3��b��#yFO���:XfTlф)v�����b��u��������x��q߶�M�1��F��]G:K���QWS+]D���ޣ�~ο����Ex�����؈����F�L&�Hİ�Op��y����9Q
�4#�>�3�����%����P 2�D��6�c��:�j�F&�����7���\6C�$��B�0�TSF�|N��eRl�܁�e�eL.'=jR�1�8**��jg��i�ڻ���g���[$o;�$8�=pn��G�c��wVG�HLsx��}3:"�7��F��a���(�S5%�eݍ�X��\�ݛ������,ÐT� ǖ<qġt~ө�(		{xM �uK^�E��HS��(`I��K���CK�|xQS�����B(Q�h���"�Ȋ�X"]F5���Q,S�K�/����<sAE�-(�2h�i�q�/�d�<�xh���H��O>�{＋��HoH\��1��Ѵb�J����Qu���	,/���f�2卍���8���b���r1�}ٱC&�?|:�Q�2��D�W�\�����`W.v��Ѐ�LX��;��".Z��Ǐ��.TVW`n[+�&�q`�n=|�4o���SF��~���Z3�]Ra���J����5<�@�<���L��o
��|��$o^2�@�����FWܦ��Qv��1�����MH�#�t���4\n(?R�י1%e��+z�[��ֱ�o�����y+��m����wl۩G�j���Z�i+楤u��.&���'*E�SkvƸ��t��Uz�����Pr����O�cL�����z��uZh�;q*���P�&'$�5[�36e4ÐT�}�b<��W0w��W��sO�)�h��S,�����gZ1�V`����׮^�����ȧ3I��<�+6���=*�� 0F�ɲ2<�أ2� �49����$>�����3L��@Rǧ�1�L:�%������X#):�w�P�D]gq��*��9���{`�^;xP�"نǔyzz�M�"h�#(�������^q��|ط_H,���=_xQp.Q������| �ׯ���M�������������`���M�鬔KB�C�]�IM���i�ҟ��q��>�b����n���3Q�Ld*'��3�����t!�0]�SOI��U��0y�P��t�Z�W��bH�"]��F,	=Y�W�<����+��g�w��m�Ap>��Ó[N������`x�eѡ9;���E&���vH�	�Δ�Т�i�CGN �&��H�QuC+�e���q�t��y�ju^���7�~/�%Ra4G�<�{�x"º'+F��{	�$2f�k�c�|�V���b��h��E�N�W�ZF����H���KF������n\��%��D�#Uue�J�^Ȧ�����]ץ;g�}�b�֭��֊��)����9N;.�0�&H��hF���Y������1�/�춹�i�<k�7�x� �S����\�t�.v��##�\]�*�Ϧ����v)P3�g��c�"���gN�@inl¬�&p����|�$zHd=��vT��ΰ�ҙ8��|�S�ם|NZ	���V�B���Lo�R/ז7N1��TvQ��I}VLp�^�
(�u̢LH����,^�������<U-���S2�P�d��R��)gt��st���8�+�e���3�%�H|�h����k��r y[ d����o�p����w�k��N�<�SS0�<�\Z�թz1*`$H2~�	�]lLH��0�-F5$N��F�*d��	8�J�xb���,Y{��>k��'�FLm�3�) ��)Y�!dL���.Ƭ�s�4��aD�Z+����FR�4��1�k���ү�M�T�GQr(B�^pF^b�JX���ʤ>v�Й{�h�=[֧�zΜ9���~�Mr�0��Z:[��hD�B�5�#�,����oF�\�ѱ	!T��3 ��H�	#uR�!"��e��u��P��㪪���q��͑a;rc���Gc�y�zd__�n��#H��mŊUh��,7K�X���L~�v7{�QȤ��Pd���U{&�^��etOD%��1���d,w��*��d��T�[ئ:�\N��'.?���l�V�8'|�*�P���d����5Xe�K����9�c�d�Ȁ�HV�����x}v���������׷�̛� ϟ�`i��k��h����ãSC�iP�kO�'�a�A�c:�[r�ʿ�rţE:e�$��@��'d������b>�@D��Y�d%C:Â��C ���UQ]��0R��TT,�v��)�kT���@9Q`袉d��#H�0�b�*H8�O�	Cɍ<[/��,��K2)�.����4�\���/RT{���������UR{�|NHJ�����L�V)6�KDL��X"!5X�TM�ZO�	c�+�/`�怀9#&������ )骩���PYS-ѭc+P��37���q��(o�Q�9�J���;�����4O�Q5�SS��]������L��1�/֘%���4�������0��uL�y|Śp�.�n�*cQdN��F��;�ߥX����:1� �2��sX����6��,��<wĥ�s���'�M�/�!Û���s��ɺ����~Z5k�߿�_���b������˗?kOO����@�k���Mc�}��@nrJ�pFV��9�2�El�5���e���P��2ba��2"��:�=Y�ea�I���Q:��J�J�x����WRr�DLU�'`�y�J(�T~~Nv�H�@_Ă+�~4A�n�ѣ���9�dx��z�4��LהugLG���D�i�/7>G�@uY�B���U��b�,xREˡ��(=�,S~�63-暱F�ȕ�P��e��r"�!H����b�d\{v�HdY���3�U�ܓ���H]e��i��(E��l��>�kk�N:9:)��e4ፇ���]R�Eb�dG��D�T�Ű_�T�qIJq��FN"�]W|Oxa�-��@��J���zu"�P�m����!\bk���K�|���S7��v�GKʮ�,�H�']:�a3Uv%"��*�K�4�3�XSTe UR"u��sܼ�0f[�	'uC ��He3B�+���]u����������~0��r���/����ó��C/�驿��j�鼈��������r����3ra[=7`
��A	dY{��P'u��t�< �Q�[H5nU.ԯ �HTX;���ڿ��(zGÔ�-j�(�9u���;-�#Fq�D@'�e4�t4��б�Iiѣn��a���*�]824L�%:$�Y�S�<�4a��?)8��	S�"\�W�\���7��z_T����^�4��\�������f��"�J $� ٫-�SD�|;��1���a�=�fӸ�yQ�$U��B?�B.-�7G����n�.�:bO�u\�;OY%�*���YT�ZE��(�����Fi��`�:�NA}tH7�������"ā\Ir$Z�p0O��/�=�R �Zf��3Ď*i�h�LHE˔��.��d�J[4%�Q�q�/nԀo�bZBp��Q;�_�n$6U�uc�+�L�)J_*���U�ȱl/C���\Ǣ��i�]��ڼ���?e��erh�pc&�~L�
�����%OG��.8�Me�V��.ϖ<S���^L��\1���,�4�ZZ��(���6�K��	҈�Ѩ�y��L�*Tl�"ex�%���`x�s۴��Ш�6|?�/�!@2%�E⨬��ipxH�3%�U�GvL�sfl�Y�$��@��y!����󘒗����2�d�G0��,�b�� ���U���#v�0}�p=R��l�`L �����<*U�e�Zp�iT!�Q4":R�h���;�6�u?�R��Ȕl���3+pM&$JohjDmm-ҩ�̹�ӑX��Dq�B�W�qc���a$�m�&$Ҕ��J�U����r�B������-I0a�C7��Ѧ
�HŎ�#^�ꓭW������|��9-*�k�UQc��]J��F�9��+�ho�g��9��E�j�&�[n8�YB�G�&��*�͔�`B,�0uR~�o���є�SU�t�}Ѳ�c��?ڰa���*Hޒ y���YS�7�HF��G{�߸҉�KW0527�1�lހ��tF4)f�9�֑��*X�2hVLZ���V����1:�HW��rT�!NX����Y�W�׿Y��R�&W"F"�m���'q8A0����\^���1U�5q��r�d�	�[.l��3��F����8�NtB
iJ,�<S8C��M�r~3#���*:-���d$TL/	h<!�D�ja��͈�Q�<�+�a��5���R��_K�g�4��u;F�l#.n�h*�n�2Z��y2u�Q�#5P��@�u��	�I�� P��kz�|f�Q�s�l50��Sl7u��)�{e� �5�%��2����ݪ��b$[d��5a�I�M����8�~MmiXV���_�SC��;��9�J��IP�|	�27�i���ӓ�3.��U�{X+�%��͓�uZ,aG+���Z��_~��=�V=��b�[ ;;w�t]>����Ы�[�����&�G����f:�Z�2�
��<��(k��D]�DRH�,���cZ�DJ ,��g4��dI�d��1���N1Ey�.RT��b��F�@Q��(T�m��\h$��9���<�xb��f�)�J�ɨ�ar��>������L-T��W#HD�"&`�9����ŧ�^�XRc8P4|aϱ��࣑���ȗ�Y~�(��������L��e�p>��Jdi*Ɨ��}@�Q���K�+FL��nS	��J �:vN���h'E�ϔ�]>,��5ei#e-W<"��jm�+�bvU�RaWQU)�E�-��.�D$���+����z���m0\��8��)�Q��X�?��Ʋ�:�;o�_�������i9$��(F4%�rHӆGF�(qIv���d[�����!ǎ�ı	���(�H�H��&E���3�]]�z����w���#m$���.���U��������|�;��)�.8�&�:j�;'2"e~�.)�E����= d�T��@F@�ոߵ�������ۖ��B!�dJ�"�o��Yu.`�[�L�2ؼx哏����w~��o���*�@���b�KO���|���Ifֹ�i٨����<`<�4/�����9��н�i�Wﶍ+wY��f�cS��>�&C۬�`�e��1�4ni�FÅՎ="�����8���\j��৊EuC(z*�gDP���u�R�Y�ڌ7k�ִ��52���R�`@�H�S�z�)��tϖm�^��s,���Zd!E8�0Ӧ⩹�@�jFK0&$2�h��+����d�%#.Pׂ��{)����$@���qe����h�;�� D�1U�CV^��e@���E����h���A��zi�����F8sP��{^.���Pll\+E�*��������Dњ����t���s�;�F��R���G�Q��1����f�4���QEߵ���@�[�&�7�m��@Q �a�d&S�����F�ˋ5�����
7������N��C�d������G�𦟻t�>�w�+�t��X�@>����~�S�����O�D���G����ڇ��4��R�'�w�,_��$k�͋�}媭]�b��Mr9�f6��#�DIH��3}M����V�ʗڷ� �"M��r�b.��� b� L������JG#���C������)��X���v��h�`��~*B�^_�~."G���
�{S,�9.JF�Ţ�5����g h�ce��L��E��%Q�_��I�<����j-N0�b��>�G�
l��5�Jqr�F��DڪDE��hZ��l�;T*�(q�U��J���w(��`<P䉚���w�\�ߺ�j�t� ��(�{�c�\�W�l����G�*z�M:z��fC��Y���P��L�6]/�9S��ᶹG�ͼ��ԧQ*ڠݲ����98�q�mY��b�;��d$A>�<�y3AQ�x�	��5��K����G�p�����vL���? �x���o~�w�����Ϟ�|�wl �l�8³Q�e��t��1)v7�5�ڦm^���.\���&T��euX`F�I�h:R� r>���`��T�r���
�BJa#������Ɔ*����k�s��r*MN �
g���L�Cq�5�(0���y
���ݘ��X8�F����n��'����Q�}�{'��s��W��et�t�Jq��Y��Q���ȡ4��#e�3Rc���tSϱ(�)��t���J5��8?�F\���[טH`O#0x���dz�ګ���8"�U��Ɉ���RM#�>D��z�ͦ����ǴI�8\�w� t~���^ڰ8�xj�0�
�QEP����)��}� ��/���y��������(��|f%2��Ć�'������g��Q�!���<й#r?����S�	��z���=���k��w����_}�����'>���ӟ���;���S�Ia�kA>R*mJq'��ݐ)�ϠP�Y��e��Xuk���uc/���V�54���|��"F4�0��y�� �L�a�(wƄ=<i#L`�>4n�j�ـzdS���/�nqL�m0�L|�xR��u�Zc1R�1�en��HF:���MH�����!R~�m4��e!Q��P=�T}S1@��J$DJ9SO�X�3�`�]Υy
��p��Ñ� ����Z���$��k�ﭦ�l���;M 	��Y�bQ�g���T(KQ(��{�c �@�H��z=�ҵA��ڰxfH��wC��,븯�#��뺒&���˻��-�?���rK^36��,%6V}&�`��8�8m�	,�|��jC�Ija��c<E�g�;rcb�*�Ǭ�zV�Ȇ��bf���gq3��$�/���\��n��M�������WH��#�����؇�/<��{mܫ��cÞ����%f� eLj�e˖�V�ض��+�\5�6,�)ҿR�J��z��2$yDU<��n)�Hi_������Ρ�;����6
U���T-^1Ve!kQFQg쯉���`�1����v�M�}r<�p���[�Ʃ�
�J��HdE´2u/b� �"��&D�Ć��i
(R���/��Q����BC����s�ݡkL�]T�E�I�8���)BD$-�N��qђob��Q�v���= ���su�$1�cT��&>�ݞ6a^�{�Ж�����^�{�ԅ6��q��1D�'6,6^��P:h��\p�$q~�J��_3���*B��hQ��T�^iӐc�74`v�f�G�Ax�-��t����ul�e��Pi��K;9���PPk(�j���U�v�x����37�v�#7n���J�W5@����_��o����y�|ػXXLl�m3�ɚ�Lb���6˗l8wOuc�v.�c��K�[�hc�j�9��V(W�v�� �08ǃ��C��9�=�!�N��н�E'x����V ��?ELn{=�d&��^��"�.��Ƀ�ɧ�&���~ws{Kǥ�Na���B"�!MJ"8�8.�3"R� ���D)�(J���hAQ��ߛ�O���>�.A�8����[ĸ#|�V�Z����$e�<Iv�3�^�У�DhF*
@��ME1�7�����hT�U��#�ǥ^j�zq������@��dQ�*�6��!��Xs q��\F�)�j  =
9��u�qO�摑�&M/ϭ�I��Sw����b��a=�S�z���ѝ};�s�&�3QYp�ʌ��)v~���"�Ret�C�-o}�Ͽ������� �]����^��g>��>�����Ű��t��g �Ĉ���,��y�u���_�y����#�~�u9�d�j�����������4�9��6p    IDAT/����ww�+qI�j3�.U0E�g���Ш.Ko�@�E�ř�,�Ɉ��x�%�IF��q���w^I�83����>����ߟxT�,�L�I��i)Q��F{F-$��BE6c�
ThI�>q>1\��B�Q���0�ZDŪYt�p��K�t<�H>�@��ϗ"'�$�ѩÑ����ңju�>	��)��!F�휦S)l$�p����IF�&��hh�wT��-��8G��Tu}v&�2
b��*ʕ?����)ɒc���!K�kP$j�L�j�?�������(<ED7��zG�z$G>�K�J,�A6ol����F���߼m�7_���eI�i�\L �si%s���ZE�,��r�F���#�}�/��͏��{��CO�D�-9�2�\,>W�ԇ�}�g?���=����X�8��,;u3�3�"��ugf�y�j��������i��I�s_0���<h,�A�k�r8� OqNl:v=�`�s+}0,ɹ�h%��G R�*�UdQ,��"r�FmƼ� 8ED@t���G˜8���#���|�AI.������=oa$BM��"�� ����&�<�������h$UD)��\d}��E>�	��;U��	N�}����v����c���q/��;�d�U���<Q��}����+�o�vB�;��t>"��2�yD���Rz��"E��0� ��UuN����7)6�$�Rd�
&���sR0
R���<(�'�hP?��6U7%�^I�'@�^�[F��7J\,ܦ���C�HR&Q ��US�d��l��������Y��m;�uӆ�Si%�W�l61��<�>�V��y>+�R�n��}�3�=��/����ҍw���[�f/�A^� ��g㵟��'����������L�����e0��V��X��ް�<b�׬\�@��FT���6��Q-�љ��}��'vrz*�p ��������eqx:�� ��5,��c���߰PH�+՚��#L|� $E �
p����3!y���c�=&���۳��C���$y�GZ�Jy��I�2�Hi)��)�)�"	���@_��/7�h��)�tYI�7�TN-��(ҬJ�"��n/���%i#Hr�R�+Uw�wE�Z �Y�L�.���,R��.U�X�1��%G�W.8٬���;��69~��s�E�.(���TE��� �z���n�;��Y
�����NW��\�=�9�s�lD�dl�Y�#���
x�d����ڔ)���l^�d%8Z��̎^|A��с�d`���4��5���d���� [X���,�߽���͵G��o�RE�:�l=������ؗ>���wOn_���,?gT�Whǃ�z�3Y�u���F�����}�}�{��V\�P�f��B[��z4E*X���y��HW���W���H��i R���H�C)"����{gg���=��*� Z���)���^�ц� q{
S�*N+"��[���~��gg�@NO�RTQPʏ!nT�=��r"S��F����M��Σ�W'Q,@��t9$;��4�J��lf =*�J�"�=E�#�����"F4��)��$�	Q�6녞�)'� T4"�O���sRH6�(x���A{t����ξ�5�.�O��D�'''��M�r�7�������x��Ó�SL �9�O��x|��TG|h�=�wx>ߠjժ�5�|�+��^�Rĝ�V�4���Fۢ�e,�Ĩ׷�ѡ\�O��lxvl���J6��bfؽ,�c+���r�G��������]w��co��S�����K �k�U�O|�|��~����3_���tl1>S��;�Fh��r�f�\M �~�����V�ܶ�/���������>���G=�rQ��&�ȕp�&�のի��G�P�{T���!R�X����u�[d *<L&2`����y�)�u�H	�ݑRV����yw�gV5�<ޣX*�;��N;:>VD��z{���� 6ě���:NdN�|����C��4	�y�(rp����g�8��b��yL��0x2�ފ�
.��NTp��w|n�i�7���v��Pr���I:A�C�Z��T�%�b�h(N��Ć�JWDa& ?΁�x�l�ֱ��h!���Z�v��m?������Y��d ��V���ۗ&���p�9�0O�c5
����ſ%?[*�E�N$��2DY����U����Øl��pг�z��vzp`'��l�>��t`ElbN���'�f 'r$[ 0.B��ɕk���k������?���6�}��ȃ�/]��������O}�?�v��Yצ �V���'�[h���b�|�v�>`W�.�� �:>@RE��e��Mn6e+�\a�=���-\��i���j��pl��L� kAM�*�6Sthi1 �GGGJ�XPQ�|�o81p4�5j�M�FG?-��}xF�3<�\������nmo
 ��q�Zs~{{�*J ,<�]���a� L�L[4�TB>�T��s|�s��b�Z��h�iUu~����Z ���wʈ��;8�dE��%�M�9q���*��b��G�1�h7S[bDQisn�L�s�?"T��$�N��{Hd�k��#e�o��=:����B����"�ȸ6?@Sm�e�*������h�AzD�Q�Qz�"ҨJ��k���!�[C�#�:�^�˨q ܁y2��;&��r��g��W��Q�rq��F�k��������mJ��d`��rf弶yE�����*_)�"_�|������x�w��W�_�~OS^!_�*�|����������W���1lh�v��Mf��\�Ya�L�2�u�l\�{�m\�����	)W�������!e�k�u.8C�1��9�*V�9�'Hvucd]v��*��xm ��ѡ��f��榋��mlhT�lz{��&> '����^�<��W+#��yϝ���׾VёW�=�ݻ�������ݶ�gS���q�%è��je)OQ�8��E.Æṷ%��x�
�w��Yk�]x�,=�q�VU����(NKw��V��F�'7!͙^)���\�5�p6ӵ��%!�z��R�3F�7(�B�Q)Z���"��{��Y�s�tz}mM ����۳g���(E��c��z�U4�#�����6$K�	�ˋ�ɺ�b�ynE�I=
ߋ�\�'z�SVp�*&��m�RP8Jt�i�gR�Jŕi9u���P6j�O�=�#H�'g-��/�V�/d���T��#+!��T?_����#�v�o�����3�l�l�t2�_��j=s�W������o�[{O�� �g9�`��~�
�5{�NǞ|��z���6/����l;w�og���G�~�$��@��U@2C���}-�r� R��9S���U)��\D���cׯ}��-k�7�	�R�VC�lY�;;;
L�&�c&M���`��9�^��h��q�ff��ƺ��� e"P*���s�TE���6lcsS� �1�?��"��4�����i�s4���L�V�b:�E�
�˿5�����P�t�������X�A%DeV�4M�͊��Ǥ��o��1�0��}C<?���@�p�� ׃��Qq�zmQ" �ZG��Ο}�i�2~E u������h��+m� wr
nvy��F�0�G����
 yޖYL��;�1�Y���܀ HE�������4��p u~�|�ו��urlw�{ƺ���dhd?r.��Dw�@Y��2ڬP�����^{�џ����j&�ʙg� ��bQ�v�z����S?���^��?e��Us+2^عpͬ�fϽر���s�̭S{�-��}�5�/�W�{���]�r�z�,�c!�)s�S�U}�m|��no����dh̜�O#�dD*�$�p+x�(���WpKi��G���n1�&-���/�N4P%UB���Bl��׿A>2N�!�Q��j����E�\p��?Q��Ԣ�AT�2�Y��8)/��XpZt>
 ������cG��ȝ�-�؂�z0T�5���yD*%�,�~M�K�f�8`Y uK< X��\�sr���cW#�
�S��t��TnM�0ҥ��uR��9�%�����VTVA�8�5��3!RڈԠ6"-��N.D?���|�R�^o������׈�D�.z�cyd��j��iEF$�� 5>�oE�I.�x��9�}`�ޝ��x�o�R�F��4�}���qf�C�|`M��]�d�����w�]���W���U�'���Z?w������y*�ħ?j��}[+��}e��a35;8��מ:�gn���q����l��}�)��������������
@:����[��y0.]��Q�yd)M�T]���!
:<�|/� ù���ĵ" ��T�UJ��z���8�+���;�,���&�C�V~�L%EKЃ�Ǐr�j�)�*���\Fӊ�:Rh�n2�Z�aŒ����OH�xL�Q�W���k�g�ن�&�tU���yh>ܡe��ʮ>�tl�R疢�Da����HQ�0HC�����it�s����HO�6I����::vyTjE��.{
��\@�R�$���_[���_�m^1	3	ȑ���s�Sy��k�R�+�
8�16'�u ����5�����3xo�9qMC�����xi�\@n4��|8ք��{�:�c�~ϊى�md��Ħ}�$�V*L,_�[��f���dK��K���k��]����4����b����N��lt�>hݴ�|�7�Ww��.��q˞|vϾ����ڢ�no���RsצV�!�O����k�,�Mc�
��9���� y�txX��b��ˍH��9x"i.��Bw����!�Aņ\e�ji��� ��T1H�^ dD�vK@I�� 1��L����̗���&ADzsf��\��k��/��]�QF�z��p<w�L3ᴝ+��+' U萷�p�|5a��s��~q��؉��-��Su"���f�1M����
�* ���kŽ 9/�^��\�ȷXҵ�����C� 	��ƽ��=�&]�"
獶��F��s�ٮ�[Ǩ�%�B��^q��k�z�V�q5z5�s�^d��<7D����D�r]'�`;��b<���#;x�E;;ܷ̬o�9�~�6��T�Y��:��Z�ʵ��v��#�s�������?��W
�������f��3���/���3��No�>�qñ�ڕvi{;�����?����^�
�����o�N;�N��g�E�ֶ�msg��Ґ�L�w����|Ŕ�X�`�$��8X,*>��k�����I��r:��c2Y��x0��D��	<y�k�>C�9�z�竼\�.��>���Qy�����,�Q)�� �&�E�,�݁"'|T�����eI3h�Ϲ�xѰ��.�&b�;yU�J�����YԵB�c�����b��(�c���Pd��b����#P�{�g�+:�­	����ԛ*8t�ffOgF:Qt�����N�k�%@��(��� #xJ�!cJ��C�c���%"6�o������^���w<?��R��#�TVE�!6rh��#	�'݁z�o�`��#[�:��2ۦg����%��Ȫ����e�t�����{��u?�������[��W����/�{'�'#���!�cwBsu`�=�%�Z���J6gO~�I��2�7����o|�U�w�3��h�Q�L3w�y&�!�i�:�w�\c�f�d,�*Ra7�u�m~΂`$�2jIڴX<D�vw������n�4�.ă�Y����+�+(Y�I2�95E*���y&d�N:��DD�����u�=��&�Y'-j��*���<�����Z����C97�@/���¥:E3ȕHՒ�fs86����ŋ:��w�0��=r|���cc�OE2q��c�T+#B_��
T\Q���|`Х_�L՛M�s�ul|�������'�ͷ��|l�%�8i3۲冐
]*%O�U���F5y5�\� ���2��X�m�Ҙ8�"�΅������#9hYv6���pV�J�sl�&�5{���uo�������V��������Wl�B�����^�o���4k}6�Y��o���N������lpڱ����&Y�|�!�������4C�L�1����scY�������X�9�&��x���&�G��u�o"d n�z�N G���:z����������L��q��H���0��6����&�\��yα �I�"�/��1#�c� P��������JT.�k�<,�$�p~|� ��{�4'I�p��&Y��۷�Q�u�]�|�>���vI?� 4U��Zp��vW�?�s��'s����V�� Ո"#��������_"+�_K[��|<���S��Up�~qL8J:�xI���J�h���Ph�5���%�L!>/
��>�~��
�7G�q���X��ejAT;u��TI����h�������بwjE�I��f�"򯅭onڃ�_o���޾z�W���c}�W�b���%�X�<��str�O���:9���/X��"��������v�wd�Ӟml]��}�]���5�/�4S�+�$*�� ���Xx�`j~sr/�abAG�M >�YK�<DepN�kx>� }�j�L�#�nU$g^�`x{���n�� _�� �2
;�L�eU4d"[^�ϗ=�)e��b��'㡢��F�3��#���3Pw:nʻ��R*��Ty9���ke�@d�c�.a�@�^ �LyY���jD��}x�N��<�s�Ȋߍ,�@cPV��bDE��"�S�&	��3��?篮�$�!���2p�4�1���Hm���;�k.�I���,<c|_j���� �7H��\?����RQH� (��1U�C�0���?�@��9�}�!����x��Я#3���kN��}f�����V��٤9���f&��N5����k�u��\��B����vw���7����#����"�߿b���G�?�t�<���ۿs�zg-+�r�m���O=c�_�c��ms�����k���k�(5;��&�A$'�@�>}��z�����
i�h�]���бinGZ���-R��R���c��t�4�k���G��/(��c�ҙ��P�9q$}�p�D���G���e�F���r|�-k��y9��ƀ��)�5�7��-Q��)�X������睓�L���*@�4Y�x��r�V�������d��}8� ��fB�£r�R
�:���� �Fʎ�'
O�W����� ��k�ӧ`��qf��z�{�~�A���>ҼR)��n����__��p�:�ԟ�twJ�&����CI��OS՝��U��h8"� r�m2���,����f�S 8��ֽ�ƤC�_�c�^�N�����U�Þp�;��X����56�m��]�/՞ڽr��͍�~�]ׯw�� ����b������-~�T*���'��!['�����Zf1�J���~O�9��ן6�E7w/XmmC776%B��7"�t{���<�9���v �NNܳ$�Is�#=��}2R0X�e}|��H(�c>GJ_��f��U㈀X,�f1�0�l�����$0������ �8'�i��-�9�`��9dH�Ls. $��%@��L���C��[��"��H'<�w`/��M�,�"-�SN����z�ξٺ,U������ER�c3�}ΕM���$�>+�� �E�U ��R+ҚyDI�R�4�0$2A��䳦�!z�#Bnr�?Ԇ����%�g6z���A��%�.3
����d il~T�㙌;����֟����f��rfҵ��β�db�hl�֩�+��gi����	���eã���֬Z_�RsmZo��\���?�����&�8�<��7����}�B!���Όc�����{�v�6������vpxlcĪ��76mm}]���dX���+UeLAqAL*,{�����<i��8�!���f���>8>d~`<m��� 4��V<X.^:�A:���/p�xM��s��2(|FLJV��*b���Ťx�%"�ஔ"e3�F�ܗi���������B�}�t�e:�DɊT!���u��7��1�>��k���0 2�Fﱢ�    IDAT�k�LED���{���U���Z���u�c��pE��G2��yVAī�:e��������* s�D��lHE�������@4��"��  @߿���{�#��#;2O�W�S6�;$d�; ���^>[2�{#��r��VU
7|>hf$ހ�Z�a�ZQ�!<�γ\�r�f�rͲ�y(�N��?\�?��{���vE��(�\,����4������yI<<BcH=_�ΝΙ�v�r�Y��j�:;���C;���<W�==M�C]*Z�R7�9�#��KN�G��&���J)g�l�Dg�Ar���y���1jZ�d��1�����e�����QV�9�����x�q|T��E2���
�1	N��Q5�s��G���d�� �H�U��fĭ�9't�����pn�~A��@�4�#=��������|�a��6��3g:�_���{"zNU�A�V4��?�U� � D8�X���^1"��r��m�(�`P��Rf�\5��F��6��W����|����+�����$ ��,����G �!�Sv��X�{���U���'�<�o.us}3@���:>s��qL��jӜc SX2k�Z+[���\гY*T�P,ˤ�9P8�c���U.~�T������}���o���+
 ���W���/d���J��0�y����rtr(N��ldf�?E���Xt:m�W�~�{�mX�ذق�����0�����](�nFJ=�|��	g�%k��/X5 �{�Da���Jn|K�̢-J�9���{TAS{���:'`�޼�ϧ
r����mv�H��j*���/m�P��S�q�he��#�`��J����o)5�f�!�V+]2q.*�."f�(\j��Ve3�ҹH��K4�8G�B<��g|~�WQ���G��6f�p�D嘿#j"� R�f�)ǥ�L�{!�漖��4-QG!�J�I"K�Q�BC)%�i๬L'���olh�1Gt�tM���vUz�H�3=c�)*�O+~��S�秨�Q	�l����i��&�69��7� ��hEԖ�)��ۥ�K��vG��3�L7g�b�6ַ,W,Yo�\8� n��a��->\mV���<x��2���D�w��o0�w�B�n��~\��V
%������|b��u�m��ά�k�L�0����Ď��b1z�L��ذ������"p�X�^q�sL�r���Sk�/&RO��vVHj���A�%�jҰZc-��=��^�	N��]��JdL�L��(���E����M���D���H`��T�4�K�C��b�qN7bp�|�H����E˃,�#͡�bB �6�B�F��:��H��׫D��� �~R�9���y]��i#�v��KB�o�l��!k��l���4�J+�s���5X�|]
�4@\WS�L�����VET22vW�~��M��/e@�'(r\w�O����'�#��R@�<R�}D�1
����'��&I7�e��y�:�R牫ꄔ��Z뾇)��3��{�B";c&{2�`H�- Љ-�L�5<���������؎�b�l;;�X�Xg��ɞ�םu�]�_��+?��_������n��2~�b �5h]��{O��P*�j���r��J9����P��[w2�n��F���Z�n����iK�C
9�a������Q���u+�֬X�Y�P�lG�B�4�Ʌ��������˞O%�,k RQ��04���p-�BɅ�c7�z`�u�B�(hD��케�ҡ�k�x=i���4�
IEpX�R�J��T�����8~��(��!���Q��xp���H"́a��9}!z;�u��[2Ec���8ؠ�b�_�7����E#x0�R��A���Gcu�02^UzxV��j@�$�6�!q]� ����6PF' �F���T~����5!� e��S���{��AF��u.7�~]� ������>?Isɣ�^~���l�
�a�[��p�P>��_G�0�ȧ�{�6�(�(*ej!sfF�Y�P�V�Y��C�6���n�tFi(���rF*f���'���{;ϕ�̳6.
��V���[y��/#6��z���_�~�Ţ���g����,�+p;�|ъ���`��[C- ���z��Zf�� �uxl��w�kc�M"�owzvptj�'��ȱkV顳c9+.J&��B����9D �^�^����.��k2J;&��$�H1���b_'������BpU�d����O���p�d�����^s2�1�!��2�A�o�B "�6R{D�|/�h#Z�o�$��圻�����V�6�6RF΋�Z d g�� a�:q"�Q��"�dTY@�?��$%5���cK?@Eg�'��l"7����h ���GKü�9�2O��3@F�V��NE��%�nSE�ĩ��ߺ�Y/܈�H�1"����yhCX�7��M#eH�i�]d�s2r�>n �1�iF���b#���e�1�j}�R��X8�5��Zݶ6�mk�!���*��Js�Sj�ee������,�}ʦyA���g 6|���l��j������o޸q�/����� �����g��/N��w�#q��eo�*�x�l�i�<�T�f����?l�hxb�r������aBp!�a=�Cfa���:C�&�gvDN�c����*5��\H�;�-z<����g9�W���� 禼ڭ�l靗ծ�ϻ]�f�uX�Id��X�Hg������I?�x!�!�1*����]`��fT86�v�I����(�)�VǞ�D*�>&��@<� AQ�,`�kB�`İ����9	��4�p3��L��YL2Y�WY���+SAG�B����YQo� ߜ�s.!���Ly���l���/������/�w���'�z����s��Y(������g�h26�ؤ4S�i��J�A�X��nG^�ѳ�2Rv��L��z�q����X�<�"r�)Avl��lԠ9JVm��䴹ִZ�b���\�j2q��KMK�F�}�����z��<W(�i���:���d�/�s�l���W���[^|��Qo�m�;�E�}p�?�uZ?Q��:"� Y��M,��$�L�¤ Y� ���cD�3��Q�o�q׆ݶ����u���mD��\�|��xj��|��z���r%���۲<N,ՆU*UV��x�yG��%��-]���h
+~����ݪ�ןu�*"���VӢT߮��g$�02��[%�Y��E�#@*F�*�H� �e.k��i�!&��<�_�Y�M�6x�H�}䃧hA;D&�,�&�N)�7U=9�H�"5��(�TQX2��*�߈jyP����	XS��k:�J�t橫��S���Β����ș�T�$��������|f^E����U*�9Bh�>�`�<"tק��Z�"���

���V�εH1��.���f�8�2��|)����)2� 6�EQ�S�-+�uA��%����=�R*�����\�Z��I��������Q����e3\o2�=�ݾ�Z����ZG�ZzZ`}f�x8a��ׯ\��_v�v��|����e^b����^��ͭv����Y����^�ą��l���Y�Hk箾�����>;ݷ���G0��VƮ?W�ngd�1��|�l�lֺX��H�:��Vߺ��U+M��صz��p���N�JI�8��0ӽ�}!�o�phG�\�\[	�����X؞1Y.�i�Ґ�X|B��|T�
"��T�˔T@�R��$Q�uRUN���ID��&���b��/:�$qI3��`�]C��W��j.����Ք0�� ֈ���&ҕ�2���&Nc��O:�iVN��G$ϳ¹E�G[��5U�y?�.�If����}�ñMm����촾����ɉ+"�������C��h�1S6=�NL�"��V�!UM���J� 2�{T��2�DQɍ�����ɠ$"T?����|?לE���%��6D@��k�ٚ���WK֨U����nx+#&@���jÇߜ��}v��ظF��W�uJ�Z�a��{��5�|�j٭��\G�)I��i֊�R����/^�����o�ĸ�<�� �F�d�������Z��S�^�� =�d5�2[,H�| �|6P�͛��pж\vl�n�2�!�T����W��صR}�F��w�v����ON%P��d�Ggf��5�����c�r���s��Պgn>�H���*���F��=d�Dnݹ#�´��;dD:�<��UD�E+�R8�����ӹ"��KC4>9��3�<��/"�h�V�}��7� �] wt�D:G*)�q�qB����y�SDD�.8���1d5 ��b��(��̒�H����d����3�FA��Y�&3���4��G����ɐ�YN;x+�yA�SV~G���b
!w +�j ~��I�I��L�_� �F������=!���e.ևn�͇s7w"� �%����I�~͝�U��<�X���j�d[ME��kZ��ǹ6���ed,�"��Ȧ�ͦ��YP���)�y�`�"��z�i��s���f r����p�po�p��������W~�ݯ���� ���;��i:?���Z9/��#J�"p��G&H	����G=y��|d����`�
f�~�l6V�{R��]M�ml[��n�y�N��C���I�������M'Y���R�i�KKb�DjE1HҌY2M ��<j���ςaR` -�#R=-�T��t���J�)~�S��?�wB��1�'.R�w����jH��3�D��-J�Ӥ;�C*`y$�ZU�T��Mқ Gx��qm��+���sN�"�R�W�'�;wH����c3�\��������3s"�U�`�Q���Zn�߻���3z�#�� �U�de�y����L9�GD��I0rB�PjI��ym�+�XU�r�V 9Ƌ��?JҀ&#�P4�;P/�'Ή����_=��10!$)�
�֨��֚�1C�RP�pH���{�ɣ��p���|�bls�9I >���g�t0�n8�q�
\�l�����cU�뵵Ӌ;��΅ͭ�{��/�X�o[y�Xԇ�{?~:������%"U
)�,Y%E���J���b�sb�αMg�=$�s1!��?:�Y;Q?�vwdc@��n��V��[o����ON�v|Զ_�e�-�����FeU�=�n N�z����u�bS� ڤ�S�V�S<K�����-�?���0�<pA1T��p�=h5m%"
�Tg���,\Ķ)yD���F����Z��x6�3�>�A�/�Ԉ,]q���$\�6L�Q�AE u@	@R���AerȖp�jo��pL٩�}DG\C@F���5�����/��.���=�=�~{*�:����<m�'Q)�%U��Rh�(΃42>��1�̘��Ɔ����&u@�~8�PO(��H�9�N򢓞��*⤙7���l�J*�HT��&㑆�mm��C\����)*����+��|�j�u�g2���g����<�ztl�,�?#s]6$�Y�f�=�ь �(��jr�Y�h|n�Bն6v>��s�Ǿ���zYz��m �wv��v��'��(���A�X�fM3�
���b��y�:�}k��`ض���g��LÝԍ�����"�1>c�|�r�+ֶl0�Y�7�;�����N�۶�w`�oݱ�lnk͍%������톴��aD�"��y�/<�@� ���3� �^HP��8�I��1��g7l���@����׵PI	�ݥh�
�6�$�y���K��MwM�#��?[�[��:RAZ�e�2���^{8��
l������V��p�#J=@_=���B��7��� ޯ�GC>�4�L|��d�P�O zt�Dq��p]�#��tmJE+�3"M�h=U�dc��T�L�AF����kQ1(�{�s'r>O؝�QD���ϝFY�k�H~���fBF�T�Q��qO�:�r����vagۮ�}�y���1#k��tea�.�����VQ�ղ~�g�ީ���l48�Zya���0��e}�
���bEc��Zi6$��Ρ�V,UU̙�X�D���f�������?_�_��w<�K_¯o@R������A�G�\�X�Y�Z�"�R�,(��2�܈�H_���Z�{d�މg���v��h��L�3|wl1�|�6m��ބɼ5�W7m�)Y��� e���l2^X�;��}�i{��[:L��r���{cc��׉B�|��7];��#	��:�b�b���~q�η;��-X ;R���΅��E��� HqTɞj0r.K<�'u`�y? �7���]\��JaDE��F5]�b�a�~p1�n���2
 ��3����/S1�� *�^
�|�����VG���N������GG
�#�}0�P�*���� �ǟrM�(#dU����0%i�63���Gz���n�E��"��m��-�7�)�ű���ϼH��� �&�L9�)J���*C��Ч\Q�ʴG*��P)R��<������|�>�|qGUl�Gރ����r'S�ظd��jJ��۷�ǘu0o�g�I�
���K����4*��l�eQO�Zݲ�����*'��-�+�|���xn�|��׶?������x��_{	�q�?/�{��?�ow:��`4xc��� t��0�,�m�P��_H>:��Nch�9~s�6�Z�j�ΑefC�{O���or�A/9��`le����y�,*�-��xV��v�J��Z{��قΗ�=�����'���*i�}���|���� �I2"A\T֝vFÙ�k��W���چF��*@�<��8�s��TեS�:�o�Ⲣ�@�S�K�"gvaUS�5d�
{J�Vn��Z�E�)�^M��v�H5:q-2t���Sq��]oq��Q�l:�xx�(R�b���4�_l���|�p�v�U^N��SD**a����|E_D�t�p~�E�9�9�s��;���$	�bp_�t}$>��A�"��!�~�� �]�}��J�+�����g��r@^�"�<�AWד���i�ψdG�d^�2����g�.��&���g#+
�~�^{��{DU�'9�d� �#M�=���c�ڦ=z�uVo�۝;z���Z�9=�ɨc�<vhH�K4iGk��r=���h]���UO�S�5��Fvv6�_�2���e�/��n�76~:�}�/���{��%�z�#H�f�=����O抹�z�n^U�|��/�, Xl�0�ؕ(��?@N�=� ��]̹�٫r������.��R�a�b��نM���v�G���l���΋J-hu��_��=��Z��K�&,�j%�I�VV�W�FԘ���n��j"��fN�E��ǜ/TǏt[c2G@��#�y��:��H�PS�;�F��{�)U�z�@��ZE�<*��B#��V$:�t2-:��AR]�"5OE#�_�K�g�/����\;��P�׆�::t�Ţ�5��7�@��\�_>+_�PTTH���H�@�I!0c�=s��+���x=i T���wc��d,�9�'� ��,o9�5�AD�]K���Lj�k��M&����ǦE�F>���M�v��C���'^���bb:�ɸg��B���	�aն7����ls�����l�^/�~��V0�l�l�.^���]�0
�׳��=[�G�͌����O������y�����C�`6ŲV�6��ذ,z�)���~���Bk<7���>��Q��w]�S/6~{"��~��Y�����C�P���G�0:f���]��1CRsj�޾u:�6�l>a��L��0~��0c(R��	�����<[�li��7�YI�!�k�ll���wۯ������vD 2:1��H���u�7��Y�E2)��Q�ع�[;�2��,@��uTxC��q�� ��(��5�j�����I������U��I�)-�UEp�����?�E +:J�9���x�,���=��X��(	�Q���]pd �l�/�)E�/��>�s�:����^p�*�%3��D"r���7�4�Z#(�<���@!�"c��{Ҩ[��S��3��B����Ȉfŷ�t�p�:uR�(�X*��e�ي/���yK"H�z}�kP.�GKv5�ԈT�YL�%�V�e�����z�.�nإ�MW��T    IDATU��S@ڊ�[��T��&�+�v��n���}�;�3�23�R'V���ҩ3UQI3��z�E�+���ik�[��Ul<A/�+k�q��fx�
lT�
ſ�޷��f¤�%@ʗ=���}�`�������j�l����3dV����cM�hhY��gݳ}�{1��lԗ���"� &���������6�V,SZS5{�-Zw��B�6<����憽�����|�~�W~ž�կ��|㺓�E
�(�5|T%��}G�-�x*��S�=�n ���x+ ��H�mq!C	`��=!�o"�ũ�D���1�!@֝����g	}��I ]��sF�!�*�]o����$!�O��@,BN�D � ca*P�������})�s�Z4W��}��qI��l�&�:�I�����HVf	�0D��HB�k�Bu:iД�qU�5�d���,�fP��c,�@-�%���yV�cZԼ6�CU������S���s6��a���\;�pї����P=##��V�/l{c���nڥ��v�e��hjf���
T�O���&X��V�����Mܟ�<�gPW�љ�����I��J��V:�NGLX[߶|�j�(2Ǿ`�I�ÅMg|/���Xd��օ�|׃o<|	��� ��������䲕&9�b���y$� (!��&�	 O��=���M�[�^�'�R���Mih���2'L_, s����Ek�����6� ~�6�I�����\��}�c��}Ⱦ��/z$���@zFY��3� �/x9r77�tn��6�� ���f��� ���T=�{t���N ��cL�JF/ojkӢ(;���Wk�PWQ� �(Υ:F�� ��F�}XM�CvP#-�|:$�HQ���,���E��KH��9�r&@�J4���!R�yH�[C_��țȈׯ����W G���Yד��"i4$�!�����t��<Z�3����`����-�lS�uD؜�g	�~�A7(�K����qJD�l,y*�N��H���gHI�*�<k\�O՜�8q�U�ce�nȁ����-{��/�=W/�C��%�	�2(�dst��|S$�|R(��y�4X�9O�؃�BA���x�r�K<{�S��<��m���T�6�\nZ�P��4ό�eDIa��v/�\�3k��_x��7?� �F��̦��e<���R)�L���:g���3��c�4��xvj�1 y�N�oZ�{,r:PyйȊ�t�s"ss��فJV(oX��i�b�:é��d��,�-����W�5�ٗ/_�O~����}Ξ{�Y=�*�h�S�p'����C���cwR��s��eyO�/�ݹ���h8��tLQI��^� $�S�3I�﯂|�� .���6Y���:�S��/��"2Itd�@��+ۛ[�I��\��_
ȅ�k,\�)J�D �w�tN����p����}'�x"�U��BJ��K�LE�U ]��Ȝ��=������D��ώ��E�ɵ zC�M����U�9�ϗZFymln��tׁ�3�H�#r\M�#����8�iV�6�jp���)�װ9�̋c,�TC������ ��:&��e��E��K����أ\���]�Z��3T��5
:�c���- �Vfj"�}[�q�"H�3�z���N�m4�*r�Ti*��x:�8�q���r0�zA9�jS�2�BE 9�e�7�^��J�r\-W~�Y����8{)@�eK�)��af�S��|kA�-_�5� ݌KUkv%�VH	[d��C~l�>�fcO'=�%G���ՆF�E�"�q&[�ɐ
s�*�Vm^��,k�'m{��-�h��g{sG�D� $����~֞}�Y���(I��R�?�H{/b8p��M۾�+�I�`�� $;fhو:q2�-]̦���4��ZRe��(Ά1��c{�;��ri|��(ƺ��5��a�!b+�ܜ "wb�,��|�����T`r��[��Rt�b~�(M�0���w�Ko��M<�7���T�M���_���29p%b�bQ�RZ�*�?x=���兏��lĈ�P����RH�bcS��K`��E���8�*w=�M*�^W�
����� 	@r��xǸb4�:���]��4�՛�2�5tͦ�3���P�ڛ_ݶ7k6�1�d(_�=�/�V���F$+zh��
P&E�F�b�vxgO���th�E+�9Jy�l6tGP(H��U�����殜�&D�̸��t��nol��@�n �R(��J��#���/���׻<����}AIT��Z#W��� 	.�#��m2�Z�!����ڨ��̓ w��l<�Ȁ��\B��a�$z�*Η,[j��iߞ��g{GG���zjwb1���:9�/}��vxx �r�"H��eY__G$�|��D�;���H��qj��&�1�Τ���"���Ф�1�$���(�7�d�XQ�����4�.�F��\t�QZ�ް.("��gV&�I) cJ�&�:�v@�鋪���禔��Jt��!�W���N�(��0+jM�����"Ј�+ r5�1=z�x�H���&C_L��/A��?����:*��?�(�p�fY,K��%�P��N@�y\��TU�堵�"�=�"�s�x�dp�Z�aӋ(S`M��1���t)F�2H�2n��F�!9S�7��\Td�-;�[�Ja�.��;�󭖵��|�i���Vd6���\�IJ���/���n8Z���m�(������C9m�m+�}R�\�~��s�(����1�+ ��sI���R�F3J	���z��"H�;�2P���Z��_m-j��K���E�G������P*�Ӭj��e� �D9f����?���?9�^��z�}�}��,ôA�<4�4�e���h�ʚ�˛��6�Z�h���6����oۓ�<o��ϫ���%� l�xPY�/���� ����ۧ�/"H��!��ȯ���jնv/��[�}q�J��ۣ�.�S�
 W#-N���֦�0�'\(I6�,(��1�P��~��g�r�NM�#g�*� �&>u{{��ET�>�,*?����)R|E�E��R$�a3��\��F�!����� s �k<=���/�= �$�ėӅ�|����`� #�U�'�#bFbM����QE��&�;9���pB��yQd� ��{Ԏ���fBQgY�I���8�t�ң����eғ�F�N16�87�\��<R�> �(�Q��;�xllq���S�f�֬�Z*��G�?�=�~�ؾ��߳a��J�f���ټ�G`3���b����\i(�d�	t���:-k��Y�H��f�r�2�,s��ǯ��bk�V��ݫ��sA��E�d�Y�κ#;k��3@����";*抿Tk��ڻ���[>�����џ��+��^B|�J�s�N%�:��TJ�� �uv�:=�B�؞{�+6wD���z�{���3"�\��v�Z�y���-�5�X���h�i�>��/�W����'͍u��������w�+_���[�n�� ��t��ww/Z�TQ�A��b$�Ǚ��{��h2�e��ɱRp�v���� ��ag�Ar7R"�Ls���H	Y�y8��ϨJ8��UpQI��!��>�����-S�u�"y��y��LQ
��od�2��W��zH�����_����x�L^ ���I�[�@���w�"�"�ǵ�6 �4��u���z�	,26"���'#~��'�K�lf���K'�2�d-y�C���(���=�B�����8W�zI��uL�=)�eP%J�Bѐ���A�Z�(D%��9����&�x�)���J�����aD�<���k2V-�����N����y�UJf�=�ek�I��4E6[�ek�4��:�g \M��\�H·r��n�N����h��3ܯJ�h±����>�\�����5�v�RoZs}�
妤>����s"I_���o�Z�w��������k^�\,nWoM~����H�T���V-���*�m#z�XpT�,3����uv�z�=�l�?���k"g+5���͝���yUg�i�Ƴ�u�v��_���xkO�#!��j:_�n�=޼���,���;Z�W/ߣ�y����
�UZV�.I9ַ6U�f���鉍&U��F-��[CQ��G�R-a�Қy��3��R���<�ϩ[�+�r�$m��;�������7$,�x_8A�3�+SN�� ~f��K���;�R���������Pj���U]ӈ|�MWP֝ڑ�(����8�D�9��۷�����/���ƴ��y��6t�͊4X���t]��=ev�B��|���s`$#^Eۉ���(Oא�T�F�8[��~GR�lƝ��0<��t`}�w	Z(���j+e���)��@��8K�t2:f`Vl���%�����H��	�0�������S�M�Vŵ���η?n;[u붏��;���fv��%���
y�
��L+4����N�1�{U�;��wzr�H�V/�z�*�t�չ^E�tri4��@�V67.Z��a�|������{��� 9�t����z�o6���=o{���ߢ��	 �[{���������lnm;1Z�eG����k�$�����Ca�}ǎ���X��|~j��MF=��[&��>��ffۻwم��[c�-r돲vx2�oړO=c=f�T�.��ͭ���,|vݣ�CUO[m=�W.�-�,*�=�,��B�msk˶vw��r�΁�FY�k�s�Cw�EP$Β ����c����Kc6�^�,G�� ��R_��mȊ��8Y�SRj5�x7Jָ߭Ҽ��Y^��ͩ2�"�s�N��\�ͅ;����)�K�����P$�s�.�aD��;_|���P�����Ըnż��hP����}�U�Dl�T��EQ%�ֽ�Ĭ�m�z��qDy7��yd=�)���_���|��s?ݳt�<�>��o�g��B�"=#��:Nru���*�;��1]��:H6���=�L� ٸ5�`Ե�|��L�^�۷���_���ʶ�s�;Hn��ڦmll�3���*Ɇ�5s�rp��,zƝ�!S{��F}+�͘��~�G�sG�C ���jlY}m�6��X}=��u���;�j�+Z�^��V2�U뿺�{����[��-��� ��ɋ�{<�}�<�\Ɇ�7�-�`n
��i���+gC��ŰG�ቍFg�A�?��l��K`ñ�(M�y�ںb���Y��c��[�7������Y[�(�k<t3�n%:Jve_������[�i�0;[=r,ҁQ�j��b�΀#�67�nkw#� i�˦�X 2��⛒�C�ǉ<�']͐Z֢k�!IT���}�Q��Yg�S�>nC��Ξ
<)�R�_;k��
�#T���s��8X���5P,3#��EX��GfD\D��܏Te� H �t˱4F59^8�J�W��<�I 7wY���H����u�y��Ω66~Gœb�e/}4���*�e�-���h� ��*������S�N�)vLP$Ů��}��q�9"�(��y2�w���A�g[��U�w>#)������p��<󌝜9ɬ��?4Y�0��u[kV�ɧ�l�{ծ^ٱ�T�Fg�g�\߲j�a�Zњ���@e���Q����@�81k��ȐI4N4M7�th�_�6FS2Y�j}Ӛ;�{�.+�7�Xn�I�ܳN��ZtG6�L��6�����G��G�E����b�(?{�~��=��\.sw<lE��j���u����������h��tbs�pzb�,�Z�N�oY�dO.�Y��A�ӳ�����}���vl<)�dZ���4��ݵ�
!�Y#�#=�/U�'p���/��o[�ӵ{��jU
��+Sϲm�l[cm]����wK,�i���� �}V��ZIIE8��;h}#��X�b&nG]H{
�S+�5�_$R����TU RTJ���k���ֱ�F}M}��*r�S� =��/88 *#�";b�H,<������"���f�#pl+�T��x�m�pf�^�R
�ƕj�;ݠ�T�F�?�	�R���#�$}w�o[��-�2N-�f� �5�J�&"i�PT�彘t�R`�Ej�B��y��s=�3�A���TEWt���b�c\c^#�k��*�M�����A�,��26v ��͛�#m$�������V3�ިˠ�g���zɶ���҅-+��͹o9!��֗��r Z0��N ���} ӳ���1���D��93|�4X,�S���-r+7 �][߸h�B�p�ǀ�ղ6�y��La�w�c�����}��������[�����{O^��v����<�����t�b��]��]�x�
Ŋ�H"���#���`rd�<B�S;9�mg�;�5+��%�̓#O�������}�0�α;{q����X"E)�����T�"�R�I\�ȑ�J9W�ʉ�تȑ+�)9R���2]�(���=������F�t��}ާѻ�8�vck�������>���>�gu�
�N�<�/�X�g��>��b|j���sph�˶��!�Re�B^�u���=Q���q��w޾a3������)ba��b(��i'�O���sv`��gtX��ݩ"M��`v�e�.�$����H])i�ah+F��ED����,��Є8|�'GT��0�Ŭi���m;[��zW > 9���sM\k��d�y/z�Ut(�ܗ� -&�m����H��$���!�+��>�ǡ�͡w��en)��Xzo�K��RN"H�a��])�8�|I��b�W�#2�&�Y~Wú4�5YW �n���@��{3��&�[��c���@bb�f='�7E���Y�zx�!��2^$^OF0 �C	��06����ɔ�$����t��Ʋu�lh�jgϜ�5���;��մ��~��Z�����4.������8�pD�B!�����c�U��ќ�=�?
+<b`���HFM.�YG�l�U�,���!�|��H븲�jss���$�>�K>���<q��|��s?�?xm�#����r��Ty��͟y2u��j�'P9:<�ӧ�lx`��������:h�N����1�.U�&LzX����լ+փ�JͶ6�5��~Tc���jQ�-Xw��J�~��޷-��{O���m� �7U��--�[}�f���jπ����ݹsOsjz����.vWd$I�"�y�c/+�"mg����g�ة�����q4& |`L��q0Z��Ҧ4;��+ޟHŘ��{���S�c���T��u9��!F��sP�Gua�����qc��I��k.x��P��]� "�Ӯ�-�+��H:�J�"������������8OI�z�Z�d������4/}NUѓ�Uo�����7�27���D�,��Y��ְ>2~�&n0�v��4���~<[*�\_D�|?dT���T���$g��q��C�yF1&0��
�漗|_�VCC2�+�K���Co{M����k6�m��h��9�縶�d���U������6�p61�M�瀃�j�\��<m~9	^�<T��;���2ghc˫� �8�r�eŜ5���5�8�Ƒ;!�>+K����𗦄��md��;�Ξ�+�Z�����}� �Y\���w��7;����*�o,���S?u®\�l��#�[ݱ��;:̨I�X�*Z��0>6l}� ���ߴ�����o��&.�s9A�N�������X�J���]�z�=�W� e���-.�[�#"��kE�u��L/J��gHR�}�C�9j�|��'_{�<��P(=�`lT���f��:�5��|�Aٞ:EH{Q'1�I$:ᳰ)dx���p�8�C��r lD" ��cD��i6��mo�:��<���]��O ��( ���6::x::���o�*/�1�QD�(�ף�ńg�ƢH�����	�½���	_.h5z�d,C��ME'U{���@����nol��ܜ���E՞+���S�ͷ�y؄��{�/�_(5�$�k�?�c u߉��~2$�rG$�3�dӦ����	���op�C�2�s�36;=��.�ܰLcˊ����|���V���N9~��zz�V� {W��,ѽ��[��L'��q(x|�.�JF�:E&��3����b    IDAT̨�О�L6g���lck�֐O���حt7��*9�������YD�shddst�������/Wǯ~$2h��l6��3O^����n�|�'3�����L?�ŅY�.� ,@ӿm�aṢ����ʖe��҂�DqG�.��+ۙ�'����u�l��"Yx���s\#�,X�NaL-#�H��"�Dĸ��b��K�c#�`ߠ�v�m���=|�TM�ࣥ�^ͧ��V�v�@�8�U��>m7��Sa�*C�:&�Ӣ��v�PJd���@.HЭ�FhC&C˦��u8�^�����y��T)�~�ϰ��6%�IEN�w�붺������_�M̩ܭH��ԴD48|�{�������Y�EpH)2�-v%\�^HѤ��r<�P�$Z���"�7U}�nx�5�'G��d��6d��h׌���R�xU���J�hkGU^XJ�+��H���0��8Z?�"�CxN��gP�j{�6??�Q ��)�O�3�y-��-�lO#�H1�8A��ED�Z���pm�O�����s�M=~��'��@2쎞�޲ԑ�8wt6m����顡>+�z胷�(1��Fe���x����ڙ�Л�\�a͡�@'��{pi�,U�:���c�s˶������ۉ�+��#��v��)/B[������\�W��ү}Z���`j�������>����lщ����P�+�C����a�Տ:���
 䐝=��U���e�<]'�6<�c'G������P�[��|�[���`�Ƒ=����P����Nm�Vזu8���~�%�lv٣GO���Ƕ�Y�B��߳P�J� #'�N��YOo��8qBe���U=pU��~ITQh�"�S�!}�iӪ`�aZ	�jz�)g����2h�.>]7�	"��l�R��C��ŅT��o��RJ�F��q���qV��T�;;��-,-��rD�a�T�������a�����BbfN "�Fx�l|ޏ{���O*����ȅ����!� �g|�S���H�eX:R�%�i�r���m�
���z0&\7���Zib�%�3�c�H&���J�1v���\ǌg��	I�6�������@�n��]2�p�8�3 ����j����oڷ_�c��Ut�$�Y��-������l��*Ւ����Gݕ�#�x����DN�9?����\�M-��mil��*�6q�4)l#�|ph��#E�+�̶������qM�0�*����u~����d��|q���������C���a�ȏ�@�s��Յ���|���疗��EK �J���?��v|�RW�v:,_鷁�a�u��)�#҃3��<�
6�{˖�H�esDQ�V)�ET]z鈔�P���Ɔ��������)����0¢+^�e`ד�Ӷ��k�b���A�^T�-� V� ��5B��q��y���+�h:�)�п�3�?��ġ�.0���	��� "�^ͣ�4t��<9)!R}�%&j�9���1Áߨ��H�:���c��J��S1"�s��ޒ#�}�Y"J����AZ*�f^m�P�G�*jJ�%yՙQ?0���v�|�u>�����^���x�0�:�I�A\~!�#'-��%r��Ą����1�Q�'�ûrfM�e,�\#�Q�ښ��8G�:��h����� ��G���tbc��zI��u@��W���F�~�?(g:y��}�+_��ڞ�)d�O�#Ͷ/��J� q����Rp
6�=e�U�����fT��@r-�=R�JS/�Q��P���9�Wzo�a;;5i�k�\��چm��I�� ?8g�Lvz�R)#[��Y�Q( ���������g���^�st���>>Ry�����'wavq��^^Y�ٮ�C��o��E|u��X��'�0��qcX��N]�FQ���u�1��˪��:_
E��vf(8huYs+؄Q$Z��Z�#���.�/����R*[�J�DEi>�aBp4�=} x��&mcsۺP):4�5s�Qq�`q����iں)B�+4��@F%X�@�[��܅G����b_�"�Wd� Au0cgG��T�w{cS�l������k�Ã�|1��X5#��Z(���ƩQ�@F$�PȌ�bz��8 U[>���{��c�c�@:f���DC���o�c�8F����*��N��x��Z�Uq���TNs�@�e�����IdCNK�7�ȁX�+z��&�W&#�3
7�l� Պʓ����E��
o[�&�N������p��x�-'H83~Z����7�Tц9�,��pԡF����������]_ņGȤ|޸�-�|R�Dֈ�g%X �)��~C#H�������ak�[����gKW<�ھ��}hC���j�k@�c���yE����S��C)�����'GO���l�K׮]s�ڟ��#5�t��OM��������;[��D`3�\�Æ��w�^�!�C�<<J��tx��v����gu�R}`���wvXwjk�f���P��j)!�s�R�i6�W���.DL=��5��(� �R*X>Ǆ����U��ڴ�6v��;3s��)��Y�7>_1F���SOm�P�E�����(Dz��d3��
�	�H�!���5˕�cN%m4����@$824lL���E��S��Ud�+�9��TBA[�X��Po��Ψ(Ν�j`h© �K�7EQ��ߚ#��NJ��@;��g�h-��t3ɑ6P���T���#xք� ���U*�Pa�B -���;Ġ�㮭�*��o�,�-�:L�kN�)5�ڶ�jh�
N%�=&i��9ÿ�>$��y0G�cȄT�N�³���n �~�����R��im�i��P�v#�ui~��<z,|��:�8D��e"A (H���vPϢ�WF;�j��=� ����v'98�Im���5s�� wv붾�k��Pj����6��M;l�gx4	ac����V�Q-��A#ʫ`�%���ԉ�ϊ�U.Wv��s��/��g��|drvv�tsv���/-����R	LackC^�H�;���H�иK8��5zf�k��GJ��M�TpŗN�Dtt�x�J0Y'�R���LӋ"�煐J��.|S��$	��	�D�e�#��\������e/�����>�~��w�x؟z����\p�����D�n���(A��a>Ũ�l8.�&����N�&zl�J�HWv�E&�:�)048��%�����,q���1��ؐ�S\�H��n�h���ܼ��Cf���8�m*ZL� �z˃��ju�Xq&(.D��H-9g`�%˖R}��t��_��m��P�-��$��M��E��E*�$��?k�療kn�=�#���ɺ�g̃uj�����������ӝ�
[-�iT���3)B�H����$�g�ң��s�]�f�-W�>wn�>
/5�}0�A�g�a��b)k�b��:1l�[k������{���	�VK�uvN��&�
y̸��F4��'n2	��Q���vw��/BU�e��SC����D�c�H��C6E���2��:Ef�;�}``�������k�����)�GwT�_��߹��2�hj�z2�����e��%���c��;ۛV��
l�i>�
Ů�ND0���o�xI�l��큧g��B���a�Ģ"���N���Ã��a��DIt���;�3�5Ŏf{�_]v5E*�5E���v��lnq�&��k�8�H�36hDt�Ǥ��Hc�gӇ� j�)�Te7�ô���cH<H�̼�4�:;D��2�8}��CZ�M��T�+U��T�!�{E��&�m�}��1�K&�a�*|�TJ/-�$������=�Q	SM$�)�����
�;Ȩ޳gxc�gI]w�f������K++i�}�:ÿ"2�g'�4�ː��l�â�)z���>��'�L"� ��)����D�U�࠺�����5����[pe��f��4 H4�q+�L3r�d@�(�|nx��"�M+�1�0�������������j�W��HԤ��,v���G���#�\[���Y�#�&$"]A��� &gHp=�#�mk�[��w`�5I�G��̚=�;��sްB�iX���S���Z���'�%]K��j!���25��S���k}}��������_\��ڻ��@�ZYynye勷'&_�CE��H�0Ib:iykcS{m4�彝�V�r?�<�	,���u�diV2�
�'�~�8���Ư��І�A
�xH�O��.T~}�_``Qu����5��H�qSԞ'O�}�5m���{R
���њ�Lj˽���p�T��)S�PD��弎{�@F!�q/�k�W�f�����^$���rs{�%�O�{GG
i.���ɓ628�ML/6�'͜<�����Uq�U��}I�DƊ2L�iZ����a�d�I�C����#�VM=?E�8Ph��y����5F��7�w�Dd�G�G?01��u���-��4t��
��pkAt�4�遬-������_Z�m��S%R$�M��m�
�'2n����>[[۰ɉI��N���G�#k�.�M=d}���/��~b]�f降!ѫ�r��bq�T�q���ö��"����9�dx�D��r�	D�!�.��>퓑�KIT3rH1��[��b�y�!A���o�5����\�&|\	��W1o�B�`p�P�.�^FԨ�>)0�|
�>t�&g@`X}NWOo�kg�O��{�Ż�����_x<�������2V��X�qT�s���e#��A'zÐ`��EtPR�B^D�4�� +RSw�wr0|����T�+Ǧb�_�-��~������#27V(��J���k����>��_�ŕe� ��zŁ�:̿�\PV�v��5��*�]Y2��{n����N��aX>�#hYo_��4�QZ8~j�5�����u���{t�C�~�7X%����e��bcuM�FQ�چ'm�n�o�\e Xt#�A�:�Zf�����
.IHq"�g^�=�jOTE+l"��'�?v��P�>��k�X�$�I��OD-��z��k�Y3��*�u�-��W���yC@g�9�8a�e��ѯj5���u�#QJ�ɘ;��X�_9g�ڮ�L=i9c�C�B���뇂j��7lkN酟v��AN$1"�::�#ڟ�2�\~���{�`���CTg�ܣbcEp2��X<�������>�?��(���w�V������K����܏��#�z�ꁞs�B40/QGH�5E"MXaO��������k��A@aQ��ZQ�"����lD�J����#��R��/��իW�g~�	��GA>m6�3��;�>�oOϖ�\ѣoZ�ÕPrJ� ��t"���LF���",6:�6R�0.�7���mZEt�ִ�q����oDg~D�(��AE��:�ò��G>��[�<��,��8Bݫ�Sq��"A渟�Ȓ��P����p���gݸ#��1v����8��Pu��)��
���G̵�coŢ�m����B��0b��o��u�M�z���Y k�т��	>��Z�O]>�^��h��e<�v��߹�D�����R���v<e�C��m��5��竸Qv��p)#٭[�VW!P, �w���g��ϵm��f�>�t?�=K�IC����v�����JI�ns3�8�aT�|I����vwk���j{��*������$SP(�)�IN���4;�I�Bf]����Y ���^�Ǐ��z	��T�u/~� ��L&�,��J���e���.5j
���*������"�e>MA�E�v�,�����yW`���O�����)=;v�Q/�E�������;y�o^�Sk>���?19���~0񅙅%YvB���Ƀ�w��"��Ξ��R.��u8#?T���7�������Ro������I��0�d(!�p�©��E�i���qM1�����.�+��A�?V�"�}"�]�=�r�݄�%Š04D�Q�>1Nۛt18�UE�G�V�����sx1vt<`�H-X���M)�`$�xߟ�~*n��Ȑ6Z��D�:�����UiO���������$D��t��B���7"7"�H/�>��C3�AWE�S*"�=t	�����<␇V�M���|O��ԏ�2�TOE�r���P�Q��?�8I�+er�)��h�-��D2z�MR�5�������|�r	�C�뱞�y1�ttu����z��%�^^^�=D���������^r���0����}ƾn��I?R?i�Cҍ5�ׯuy��=~�XFQ'��Pu&Ԯv�����'�K��ZU�P��U�.hE>$	�Jݾ����r������L�иph�	i3�Y�D�|!�cG���Cǲ�.�2[uzP>������׾�'[/�H���򩉉�|��ݿɳ㓰EBv0+�G�q	KJ|�ef��G���J�I-�������#���@ZTy�����/��IJHD��<UX!���+�xUS��x�-���uÒ�**QE�O�SR �K�@Hq��O�I���k��02j�v�W�����us�6�5	^)�"<���=���KW.*����yQ(�}�Xs���������=���sa���g(��L_փC.J
%��#�4s$e�{�G�NĎ^�p���M}V�@۠d��k��q:��ۭ�	j`?�g�J�߇N�r�u��] ����k;���6�@ݣ�旗lNo�n��Ƀ�8�\�F��a뛈�X�ܣQߠ$s���9�S
�1�����V+���q�ӊ�x�AR��w1��?�1==k���3Z5��{��EDF<x�އ�5��1���KN��s�G��o��s�����!��0t(G�@N��`�B�N7Ӛs��(��cҎu6�_u-&�;}�Xi���������޾�������>��'5���|���go߽��[��~lck�/:)]����/S'AFEnԥ��T�Q"�N�q�U6wxĈ"� ��H�W��X�8U�1�`�`1N����AGZ鑥�IA��Yw�l�ϟWqfeu�޾��--��o�ony�oJuhv���C6�@o�W�i�(��E0FDb?�EI�![�^y�D�y$��F�"�p܄��w�%k��C��tznZʥK��A�0\�J�T��`�Z�\�Tث"�N���;��g7v��yB�l�mT��e��i�B7��p���U;�q)?^˵�	�A�%"J���V�'
=
:��̨G�S���/8���S�)]��GĽD1I\��;����zq�D�K�Z���-a��ż�v\�P�Ø�f���Ԟ'��:�0�0�'��	���2�}B��~-{�K�y[��u`�s�"�3�(Ѡ�{�ӣ�599)c�5�H
��W�9��_獂�X';6*��N�"rI���K����	n*��>*����,!+�(~��]E`����D��D�׽!'6�E�4�����ڀr�u��s~�s�����5�ߚ����;7~��䃳p�xp>��HȫjH���  G�X�p*p�ljR�X@�R�0���4�}C�B�-6��K�+�8�,5q��XM�B`C�G��14:b�?������������[][Wj���⃥�)al���+ �a��0B@�	��Q���~J���}#���;����Q�T���i�zͶ�V�3�RQ��*u{PT���YG�� �Ch��k:4������s�^��IL�	�`�hH��R��h��E6?uT�'Ġų�5�m�;KZQ(�!a�A�qCI:��|C�8*�<Gp�MΓhM�q�ڊ��D1&]�*۝r�1G;N(����k�k.�娈Np0K+�673-ܑ2)i�*�@�G�k4��o��|?` �Y��{��G�9��;�.U��Td_���˥�3O&g���@JήPl���ѣ^k:�C%E��`�qte7�@i�伺��L���SV��#Ux��b���c�T�����):���Fp�B��č���Zm��X�A;BSzd ���ܯ�wN���������^}�O�~��#�f���wo��w���<����@:m��A�ԇ�«�<�S��s    IDAT�1�v]PQKj�����=��\rIi�ȴ�οr	}���mn��I��H	�D"���K�<P�3�<c/������w�|[�~�V?E{V�c�
�
X��{��C�~��k�:�p��x8G
�S�u��;C�u>���VZ_�f����v��Wﱹ�#��Z�ȵ�$|h2�5�0+�F�k�0��Khq�Kb:���]'u�EFd�j�j���U�DP��ȁh몡N�� �C�h�
���Q���ob� ���Uq���Ҹ"�JY������rR��(�aރ���$�l266&L�Huuyɦ�[mwۺ� H����Ξ��o*���B���9����b�V��ۈ�
*RJ�IJ)cݡ��k�VN�cuY�<�9�!�Lk�����7n��F�@i�����T�R'�	�E�z���ո ���#��!���"��z�$1��1�2��J�S�.v"�3����
�IC���;.���O�5<د�����Z�T�sv���ׯ]�gI]$��m 頹����7n��/���v�̠��TSj���{>��}܁�&g�ˁ�t�b0��[\�$���6Rz�}h������̔�kP�ҥ��@�N�Ufqc����!z���U-������1Y<"��NO	��~��z���A�G�x��M��"t��[t��pR"6$R�����%;�߳�RA�@��C�,c�"���ܼ"�F��fS�Z�T�Z�bI���ދ/����Ɖ�M�tb��Â�@dj>�Rp���(��#)�h
��D����<p�|O���1�E,�	�(���8�A�t�����x��Ζ�wPJ�Pݒ-�p���y�=0iN�5��Cw��)+W{t?ˋ��������2�9[]۴p���hR��t���A�T�bR�dE��������@�QT�6�eҬn��pR(�0��Z8�ȳ	V�����gǌq��MD��S��!N~�<����%Z����&1�:��+-��5ʁ����oچ�y��).7���E_�T���cgό�N��������S���+��'_z��s�ׇ6���������wo��+k[ۊ�A���W)��&	-"&m8fOh.ESx]X}�i�H'P�T�����
X�~Q�L�:h@�6"�Py&�fQ�{�e��#t��\�b�.]�^��{��"6�p@�=z����#��!d{��P����%��)RT��孓�3?0V`�T��{��qM��G�x5=��U��-a[�wI�k}����FR���t�ҌhY�r�����`�BW��XUԺ�����E�J�bӣ��)�^Dcq "����}VK+�bmP�aצo�?���.<U�9)�8����;%0�@XXہ˄2�?~�ϼ��8904����J����].i>��q\�;�B��݂�)Q
c���it22�t�9����"ƀdRĈ�Q&�d�5��魟��Cw���pV�뭷$����hؒ�p�:cT�+Z����OJ��J�+.)*�G]cocn��;�����4Q3���<ed۲���oL⅛�~�>S��@�jc�N�� Ё�s!���x����;�ϯ��ڿPX�C��޻w~���|���u 5F5�1������J��>�B�案�νJD`���D^�X���a�\c?������3�Jrp𒡷�d��y+��B�A��p H��>}jSӳz
~%��m`���1WJ)��1%������i�w�!�	�%�k�S{�=���rI�G���5hq�����1���>�5�mvv^�0��=F��(d��Y@��9�P�蟸dJ�KT2�Fu�3��TF�<�&E�c������K���q@e �������K�QS��X#f����8�W�����9�G�:��F���t4��Ԣ�{E=��LK�,^�ϔ����r��y;}f��{{liy��=� � \KĔi�=H
��!g���z��'j?e�i
�j+��?�(�i�G�89��`����#J�H�݇��s��S�Nm��]���u�xּgLrgyD7���2��k�X��"�~:�3�%zU�[�p&^�qU�x��~�km��R�3��$����`��+��W����'�B�KgN���������d2��^c����ׯ�p��_����rECw�R����ǡ_��n�Ԛz���p>�
����p
_H%�
<7���A�v�"&6:p�&~�*�ݺ�$�zp���̕eX)άml�qHc\5c8y�^pͭ
{R���;~P필���m���CQK�p����}��aD>y~^�+?�c��N%Uٹ�Emv��C��)N��3�����{�D"d�S��1�O֥�1�Œ��׏s�k@�n!�;����E���k����"��fҩT-��
T�$���L��IM*%��5"H7b�e	o���U-��=�a���>I�ա�P��k�hׯ_��@݉��V�������s���L=�C�O����dV{{�-͘�ݭm[��u�x�1��n7���� �
��UEN�JM~�� �ϸ^�n8G�VD�D����<��A]NW�^9|���c�9�1(I��3:mNt*����8����2nO	��hZ�?�BRu
���
�>$���36��ok�˶47kK�,��������'�'�/�}�A���|�'O��u��߹����]�9�C��K�=EI�H�-�����^#>�� ^#E�M�E"�����E�("R<#Ə6���z���3���w��i����b�~�6��,R�J��⨴�!��l� ���hϣ���f�C�}J�Hy�9;=v�F�G�茡C��������3g����5I#�V���-,-�8��Z)=N4u�0��i4^R��rsEƑ(V��E$t��リ���9�mc{�667ݰ��t�d�j���\�xF�М���X�Σv�<�r�� ��}�������-��q��ӫ���)Uu��=` ��H����(Ľ��g����-��QoH��҅F4����)41'rC�G����k6=�D.��0��+�N*>���@�,*"�V�s�S��C�7����%�u@BjC;�}.݄�X��Q�t�5o7�(���%�n��J�^H8�*�"�+AI	��Z��]�S�J�#�Is�����TJ�Xd`�Hj����<1"���h󳶱�,�h��R�ѕ�����Sg�4#?��|��y������7߹�1U�3``=�T�SG��3\T���zy�sޤ)�R7�5������H`BJ�y�n\�*o��q #}@�#���S6���_̜����̈H������Zy@:X���T?����N�	o�{:`}��Ǎ���k��@)�A�<_h�J�h�J�(Llh�/<o��mec�f��lzaN���J��ѫ8�Wb'�i���F�ӷ[��@�W�����vP>����HhqT�pҰ4�2R�H��f:���<��1L��A��.(��h��q)���� ׯ�uȎZ
E5
>��\�̆s�(��%Ė��}��~�&$�f��- x�;�V���>��������oܲ��!�۫���mml��`����aS�)��٨�"���[RJ���R@:a9�Ni5cr1��=e|D*�(r�I�`ށ��r��ϜUI���#���H�(��1Y'7�a ��Ҥ�����W���\�-�b+�L�MQ̉`��J�O�������^V2�a ��6P�ة�V�Z���AS���庲;��\��Kϼ�K׮]sNa�Ǉ7���/~����o^!C��]V�j��ȡ$�F��A���R9�r�x~>x82l�U�'�9�ikHT����#<���j\,��`�n�|�@�ɀ�q��1�(���P���w��"����^�'�DR?��l5���F�a�<����Ο���c�S��������Ǣ�Pm'��_f6��-�.ؐ$��1"D���;Z��ct�W"!DgT2�v{}��W�"���b�M��L������ad<*�7]2AF�H8�Վ�aJ� �Ji���+��⇻�C�h3/HQ��E"<s�y��� ʥ+$�"��$��]IUs/�PD�y��>]�5wgz`�{ެP,�瞳�S'e�����
Œ�G�y�)F�l�o�vw�l�@1�G{6�=F���ڛ;��j?x��bE�I��
L~�"��T��@RgT�/^�(þ4������q�Q8���׺�b��̩�D�����Wʜ4�1]���w� R�Gd]Q��L�=k+�lyzwda�:Dlry���Z����[]�W<][`��ϟ�ߟ���G~�Gf>rykv��o]��_�}!/��b���+s�9:"�&1su��t%�O6@���GuQ8Gjy#r�}1L|0?%ں�iR
U��T�����t����iGv���8O�N���|�)�?p�ک�ǖ|&
7ǝ�@3�G�gyA����BD�)6���а]|�]<Ϊ��풾��*:!�=i˫K���l3s�����F��|3S����O�T=��G*�3Ҭ�fS�O���42E�Sޛ�1�Og�mjjZ�!<$����h���-@���)H� i]CG�J�%�fB��:I��8�<a�uN��������5O��G��.���'�ׄp�B���X��"�K��(M��whi�( z�_z�y;s�����u�_\�г����W$N%��ᓇ�U��"0��=�q��a �)@�|��R$�~t���"#�B`����L���S���t��;�� �L�3�w���>�|ƌ�Gix]R�'��
�Jb��}R�n7l����C#�LpC�W�CO4���~���bdG"��U��s�A�O?���%E���=eR�O���/~�g>��������� oL��+�o���oݝ8Y��|�[�X��$~�<A������ �O��4e4���1>�2��O�+R�tυ/$�?�Wz�d�������%�'���eW����---������Y�b�;c�i"]z��o6axi�t\ץ	x	�$Eiut���2$�ۆob1Rlt���E"K����bьƁ�.���ڊ��׶6u��CsE����P�fSk���UF�8FH��?<���+W%��M��d�Ƹ�=h6me}�?�n#	��{eS�jD6�7�^#	�����0��X��\��ȍ�E�Z�)F�Å��#E�s0�^dp�#������h߀T�ٖ[��!'��5xE���9��iIGQ�C���-���?�	9�����tfVb0���I���%FJ��z~[�Y�M���<��j+��yr���vq<|���F��8��1������y:m���뤂�Ul�&_���+2L��
{�2�S#�h��s��="�y/:�]��{0�]YV���y�@�L���)�����=�<.���pU�>=�����UE�hccc_}�����O��_���#�7�f��ͻ���Ç}��W������uy+Y|h�f���BEh)��#�h0�Q(z���,0��$��>~�#�Jy,�R�:��9�^�}6��/�`;ۻ67?k�K+�|T-���}�"#3��f}�!
���^��D�v{�������1!e�}�S�>��g�N���W.+
�:�/��hm{�& ��m;�=Ov�N�8s��2��h��Z>J%z�h�;���t�@�""`t�I�I�%���_z�s�K���c������=iMn����#U�i�Y�ŗl�r�g��6r}p�䔈p�y���Nӥ"L,]��;K�Y��>V�An������"�U,��t��+3��+/q
�z(>F��"@����)�@3gϟ�j��S{�� ���S��&T�jc}��ܹ�D��Ҭ}��1z7��H#C��YAH�<�{�ȍ 7 %�8t��E����l��&�����=�쳒@����F@���TdI/yZ����S��t������P ��Ŕ�������171�3C#L���3�8_|����q�z3Ȣg?����{��g5gsu�6W�m~n�L
��������}�����>Ry������s���������6`��+綑T��d)��y������*���)~GJ����Z^W��A`�@� �HC�<�i:�)��@�����"!<<i6�]O��]
�4)Ĵ�0~lT��Њ��8�-��ш�d��Ұ�Ό*�����ܙ�J	��7,�a�[�uu�����{8��m�CZs"��΁فmʰ�g>cX��EWfA,�(A#(�e:�k )�$#��M;����������S3�9h�(6��^i#��F�H�t�� ����8y^�/ʘ�JGV�H*�Ɛ(]wǥ�R ߒ�����4���;�u�o���G�27���K�����;~ϔ���:p�v~�n��x��.\�(��=t��]�By��]�7����[ʈ�+ ����J�j�[{�:	b`|�1�!���R�I?.Z�Sl�{���w�`0�/����]�$z���-�A;kE�D�	W���B���[Y��I���yRtჳ��H�j����d��982���3�C�MR�D%Jc�]'��`�_�j�Æ�l����-��kuOoy��ŋ���3��>���ȷ��z�N>��&&��++�-��V&Eq��VҜ��X���f1CT�6'bp�H�[�W"�b�c���\�Ta4�ƅ1��,%�o�^,�����S����u��9,\_�����N�^j�\(��q؃7�A�z�TT��w/u�+�UT����A�=}�.�;+p��tox`@d���ݘ����OQ�����+�� ��WZ� m&�!��uJ�%_Цf��m���2�D���e�0�SOgmb��#�G��Ҹ�q
�dI�':����v��^Rzpae��C�����S�F3��0�,����A�����H���%)����&eV������Սu{��i:|����Qƺ� Ҭ�#�jfD�	�ⱱ����K�@��K|�b��Ј�tff�&�O�@�瓊�9I]gd+��0ah�?Q�=M*���1��gU��=���}�W��W���Ԕ-/.��
}��Җ�����Z�q�!w�_̀
@XF�9��~�V��Vh��P<��`鰊���$��:�>wEb";붺8g+��6jvf����g.��+_���6��0ȷ���ޙ��w'|~��P�ձe�j�k���,���g�$8ᩢUP�%�ű�<�hS$b)�$�+����__���w���a3T�R��u\8w�^{�5{���E�O'�P
�i�צM�QDt�!=r	t<\��f"�UH�.QphG݅�� �JJ`���K��矽bU��+k�p��T���u��o����er]�.�*R��1<a7	��=E���#�06b��q��fSFQmk��",v�˕[4!�p�����f�` ��C�"�������y�
ÛIDD���!�=��%x���U^��IM=���Q�g���פ�P��Wm{}�vq����*U�W�(K�����5N�Nm_�1ׇb���Nj5ɸ�_ͺ��CU����%{�7dt����k}����G���I���?�t��l"C���U�I��0�Oa ��ѩ��<ؐ/���Z������R�0��[����'G�g��A��0��<�@F�}��c�F`��7E��u	z|38�W(�@����?����g/[)��S\�����E�s�O?�������7��ѣ��}�O��#�o��Gw���q�n	J�H�!�X��6s��$���V��Ns1��=��#D�,J��TEO�Ǌ@�j�>�\A��1���(O���}͞<y���s~����1�����$��?U��Q�=�C��_�{D��O1�=��k,��9U|�#h^~�y;9<b�ڞ���B��6���쬽u�

�L��:����V�Y��h�VW ]��$� sY)���T�љ���k O����J���'T��N�j:���TD����sE)mcq�Y�j��HD�Β`������\��y1�}�B*Zml�����nl��IC�opHrf44`�h�H��i�� ����$/�    IDAT�ϳ �e���"ǫW����'4��֭[��o~S����rv~�M>P�l1��;=��I�8�%)�e@JQ��aV�B�#�K���{2�#�(5�(Hb$ٗa# ���B��jL-,0�Ĥ 9@ƿ�z���č���H����t��qo<�1��IRo :j��]PK�}鞸g�.�矻bC�}vX߳���m�r�Ύ�|�ҥK�3�>����@�Z\�u��/߸u����=�U��q�	��x�Q��`q.z0݀�G��N<����Ʉ1���(B�v<+��I�!�Ͱ��9g�s�t�����H���g|DxOZ�k���gu��j�M��;I�X�4)� RPwB��Bv_�h0Z�B���΍�����jc'N�4A��N����=9iw<���I����IA�>ZN�p�$_F$�������t���lG�3��?$_;���q ��f�>xl7'����e��o��y3^�	�#J��UQ{����Gt�ĳ�0a CB+�`+%U|V�E�B�XrV�-D�Zv	� E�5|U
[T���c4�͛7E[r�ݥ�sɬ	gL�p�{	�AX�+�/ڧ^�a���W��K_��d�FFN�wg������b�BN(���&���U����L��#S ��_�~j�kیg^�[;��;�C>ME�6�Zʀ R�����T��:�g�����QTc��9j�E���0����ʇ���0���=��e��Fb<y�Ж��l����{�.���g~�/���$�޹~�޸}�s���$�1}��2P� ˍ�Ј���d�B�%��a�b�Z�I�RjF�H!�74n�P���O�u�\Qg�P��5T ?��뚿��o�7��H�5DlwW�R���oƦ��f��hz����7�{|צ�����[)�Uy��%;5zB�������b�'�����&�1,MP�M!7����8ئ RS�X��/�`�_�_���b`�IU�]9O��K���@��j�b׏����v��-�]\6��"��թT۱;�����]85��{� �6`D6��H�镚�-L2M�d?h6>"�4bh��ם�#�Q�݃hU�.MK$�>!�r����:G��:E�f�Q��5~($G�6����-Y��_xQ���?�ïk����19��y`"Π�E$dnAQ�\I��-e,�5Eo��(~�gf���YN-})h������uNN)i��!����V�2���@�w�<h�bS�������A#�N[��0���Б:����Ɨ�n�$�sT���ٳ��L=����%�ޙ����¹��x�b�#7�7ff�߹q��7n��4�f��,.�A�"'1I���@֙s�ar����G��u�M����cl��EtU0E,�s[��&T��GUgϞ��}�c2���o)���VB�ڽ=L�r�B�������*:$< B.E�#�5��Nd[�Yo�"	�����m��)�3��Εm��8�x��8����0\]BJ��@j�RJ�qLj����6��T�B���q9;6���1�P%@ �@��xԴ�{��c 1�ip
�Ө|]�Rc(����?�趈�2�(H#�����*�J[�B������
:EW'*�VF��z�,sL0��b;vr\��ޝ{¢E�)$][@3���5�nnȱ����&r=���^Rfr��m��w�#��f~~�nݽ�2�aC�%
M���a �Ȱ��6bO+�M-��������Үhv���g"H:�B�.ddf��Ѣ���M�2��P�������A�A�b�����bj;V�n$�w���1�Zۚ2�(qt��3�cvᙳV_~:%&�a��`tt�o�<�[׮]c4��||(�����}��oޝx���O!$��	Y1݌��{��+�N����i��c�����x@!�NQj���4"#u�MўR�0��$|�J4���߷{���9?�CH�"�op��9Α����;�JP�UaH�e̓[8�
#��HA�E���V{ڥsgE�)$b4F���{�x~Ѷk{����
iU���=P�GJ���H\�3��D��kk2(@C}�2��RA;�h I��NL��7������%���3�̞N9uE0�=���F}(p�����@��e4��"��@*O�0 ���R!*W��Ul ~����A�@ԭ�2������w�w����"�f;�%�
~��]E���5����龞{酗E�&����-��V����΍�Jc�.�5���'��p >
�X`���� �r�5��))v#*_�D������V�A\G�`g D��^ԉk�{~�Ք�ga��q�,�u���F��J�Z.C/4�����6<<h�C�V�e�g�wk��J�O���;?��?���~|(yca�o��w���]4��M=���� 1��?�!�AV0�y}��ƍtUHZ�4�����?���8V�QT�ҡ0�a ���� b��<���J}޽q]R��֊D��D��c4!��4�v�'_��h�a�d� �W�@�=h�RW��s���66z�t�Ό�NS��旖��Ą=�_�]68�?m4�a ����R�M�v�l!kT|1���� A��)�V��+�"H�4��n:����-Yd.K���Qt���W:�ѭ�e���ҵ�����>J3u�d��#�����=HD��A��g��kO�1�A��M�>G����c'FF5=Q�۷�
�ޡ��9�kR��sp ��E�Ԭ���@_�]8��]�|Y��ۿ�;�z�olm�@r/����[���F�h7�3h�@�}�ጂ{A�<��Ĺ�^M�8N���A�Y�f��C���B���3ela45������"K?�mXZ@4ƽE�$�ڪ��*�J�x�P$C���UGZ��[�2���+�B�0��R�	k����G��|��_�����*��� -���D�y����"��P_ϛ8V���s{���)@x y��p�4%y� �j�YtD3���/���(>�Lz:��	�r�f�'�d��;���ȵ�+WS&���fbT��Rk�hR�k0�r����s9�x��=w����u�0�|<e7�M��ʊ*ƈ<�
E��*�ul)F��H����C���^�X��ƥ8D�-���#�x��+i0��;y��C{��ME��J�erE�15�Z:�>�!�|��L�#z��Ύ�N:E���[C��g�#< %�4q�6Bֽ��W���*ܢ�`��sHCD�Q��s��\ֆ����T����4[���)�DWd�pumMn��FXo��L�þ�p����W���VWT8X]߰�ׯk�}����(^�z��d��ρ���7A�qF�RÄ�_�B�<a}}��|~�ޞ`��(}�Ց�蜧6�V��Ɓ�sų�,2�H�ym�d��y�{�z:c�H˗�&�H��3I$�jd�Z���A��AS ���]�����㧮��J�ߏ�[���;׿������� {�h��ϒ�B;`+�d:1���8�1"
O�������J4��?�ޣˣ�P>��G�'cJ�(H6���ž�����'���hP.b#s] �J3HQ�G�n�&8
<r�yȧ�ḿc;�V���2H�'mH(7�ȮƁ={�={���t��oݹet�0�����~S�(E��|c�&
y�����z�yi����5K�׍A�H�W-�w��[��'#B�ă�� 1��R�2]^,�t��Z�ʧN!��L�uA�C&"�8����$vDD#�[�}�@zD���%'*�T|�=�G���b"5��z$�p�yT�d'O��XAN<��b�j�4�L����r��Jvˉ���I�3J�_~�{�ա~�T̷�}G�K�VP���AY)R
b>cDi��F:�n � �8:��FhD	�Q,�{px�0���c��Gu�q�g�{�1�5D����9>G�^�!NEZ�/~&�!|=�Z@?��z��{�5`�#C�6Ї�iqi���������իW?{�H"��'&~�o��kSs���Gh���������i�r�0'���B�9T�Sca�ۈL��C��lھ�~����Ek�
�ؘ�X��E��7�aS�Oe �V�Je;U��.���q����E�G�"
��xI�Rå���Yȁ�?(Q��-c�p��0����+ϩ��� E���-�5q�OO�n��a��)��$�FJ'��28&,ң�l�a�J1�f$����kPD�@V�%Ž��u+�h��0�;���M��y�JS��Bz+�8�@)�~���f�K2�Yo>�Y�a��CY&����v�lo=�;3r�.W���u]�Gȏq�"Q�0�Օ%E�T�1JT��C?�7�zǪ}�j�D���i���,^�Z�V��a�2GR�����v�'>�I�5�f��/��7�#���(��G�{�=m���'*�H؝eb�DQ$�L�8�H�J�H� �~l�b;�ێ�GZ�n��#���8j���kz��~�6���*L�8�\G@/�<�)�=Q�o�#�0�V��S���ުu���C��_�80��/^���A~�w��s�֯�,,����Aa��1�F�l��{�B��xs�/i��I�;$��3��M�H)|{د�$uh�}o�?��a������h4��T��g�(���ܳ��?~]i2��"r���9�����Wܹ� ۉ 1������6��i&�2@�#C/��;�����h�+Ͽ(r�������=|�Ж�<�`�\���ޠ��4�!���<�~*j��5��"ⴹ���l��� u,5�d������7���Ҳuu�ٙ�f�����!���` ]� ��P�L�� v�����T�H����c���&�*�����/�5�?
:�D2�{D��H#I�1�����-��J�#�##�[����?~�J�^H���GȢ��!Xk�*�i���i�==6�? u�W^yU{��o~K$���M5"����p\��h�ù�p&8'��czLo�N��H=�
O`�к�@��|��������:��3�a8�0��.�>��8�4n(Շ'���q�Z�O��S?���P&��ԛ~�hC�;�BR�?jD���>�N��GF�Z_g�_}��4W�-�� �����[�&yvqi��~�4���'[HRK��Te�4�-��6��H�O;֋k��-�@�ydF�
4�$*I��#e�l�1��'l���a{���W^���
5[�;j?�=�t�gU�wh+C�+QAgC�)];:ҡ��HBD��9��y�N7�|��G�G�vp`����]�p�{mg�n��G_���U
�#�e��"������&��������0�2��]�"�j,�� �7��y�Bty$`DdqL�a�n޹ko�x�{d�8l9ʤ��xtdDe�=��@F�0�y�*:$*�jO��v��]oU$�����].[�ح��(�_ΤÄ��:Ԧ�7�Ԃ�����>[��76�UкS��|��ST���km2�����S��]�|Y�����J���ʲ=�y�PG�+�d�f�$Y�����É��@z괚0hHE�I�U�!I�R�HVpdP4JDv�+$#�e�$z�N�=��gE@��Ge1�Dp��k��Kڟ�E�)Ho7�(��gOa��x��|Vm�S�ld�\zr�䩟�����ﷁ���O�����K,�6�SjL�[�y	�� �p� d�X|W6�4������t���U�������_{�+�ڒ���=�@�?Ky{⮞�#��}��J�i�9Rޠ��x/�P��3����3�~�= <���v^j��:�5���P~���\����ַ������.Z�ܭ(�9�	l�(Hp��p��P�W���,	�44��G6�%c(*�zS\L*�P�Z���PCk5��q�=]X��b����1�rP�+�t����j��v��{S��4� B��������I�覈VUp]��ƺ���;�Z���o�Kz���� ��[VWԳ��<Tv���V_��75���2V�ۛ�A��9{*p�=Eɜ(�T�Fo�.�?o��l_��mj� ���%[]]��ǘ�0�����H ����I�[A�{�41��#��
�N�״���X�^xA��`��]����a��r��&G�-kLt��9�|�ngH�Mʭ��C:���f 1�QI���ОIjK��e��@k(JY��c_o�ʥ�3��?;�����W�ͮ�o|�߻y��=��\	�^�t $���6�1MWK��Q�����U�o2B�+������� �1�:��J���&�;p��l�}� ���^�l��{�g����q��rD A�F\�a�m*DY���3T�W�.�mZ�ؤ�Z�Hb�E�dS��v(r�e�;����j�.^�q~e����}YkP�l�(cG��up�a��s:�-���M�LD���qFeP�ps�B�z�+�d�bVjsS��zRvpxd7oݱo��-�oZW�[��(Sj��ѿ¼R�B�,��2�m�SD)rPm�=`�<kE������xD�?���~�f�K�����/��V:�<�R�[cJ!��|1����)�������Z}獷lcsW��1Z�D���(�/8�z��F9i�ʅ��7��{����ʊ�{��#sxO�
�6	�s��=��q��|%�����d�)�x�r��b�J�KI^��x���������TzR�?3�,|0�@�D�2��m��Q{P�Ϩ�$v�>`���^�%�a���O0X�1F���CkT%� LX��Xbr CW�t����T������:��s��_��a��?}Z���4���ϯ�md� *..��B)��Rc��|��-�����"�T�}���>P�K��%6�"��3���+�MT!Tp��$*5�e��I��O�R�,
���i�9��CAGƭ��C�3�1�DƑ:��nO�5]*zI�D�7��$��>�V)��՗>��^"�����?���7�#���4:R�0Fa(�Y��M�����1�U*�fYfvwvYo�[�2�CR��>8-䝻���}Ӗ��P�&��:��N�W�<����2,m)���h�K�$�j?�X"<Ş�>S�?��C�8�U'\���҂շw�F���@��MT{{%rK�L���A���Z���%��5����o�����m�M!F|htfǸ�u�uE�r�Zo�W���jBx�;o���ť%E�t����=�
B��m���)�� ��k �Y�t�RS�=��FRm:��H�*��h6�*�%2EL�q#yW��ȳd�q}=U�����.�4�]�n�Za9����2�B�� �@�����K�7�:J��Pm��#��-W{�3#��=74���Ν�q�/f�[��Wo߻��&N����NW���A�@�pIq�ѥq�H��(
V.;����79��
�KF��"�+P�Ѳm��xm`"�0`Ɛ^�o^w�g��ի���@�@�1�T5>��-T��lj�J��>�E���r����A=��S��s�Ђ.A���ǀ"v����O��k� �$�?��w���X��ݚ$�0�j)L�?Q�¸��w�֕~åD��)�H}��*�
Z�U|ɫ��Ǹ�{�о���6��bD��&� A7J�[�-EA`�J�#���5����"�'Rc�/K%���4>�'r�ޅ"a�$0�á��vg}S��Qĥ��r��"p������-.J�0>~�:3]v��[\Z�z�udm�`_������ �N�ڶ�2-�5;9�&���I�ܟ����3R�0������T���&�����l�C�,`���-h(,ll~�����@�)g�Z�=�"e܁	(*2&���ƾ�wo��Ś#z�D6�g�5#���J"�����r�{����b~H^ы=���9�'v.c�GF4���\��Oz��������A}��zn?z��<����FW`D!5E�8 1:�l�-��Xv�$��/�5��@h̍xgVs�V�ΧH�����a3���Xp�x/���1�/(+��_U�Q�ȱD�I�RX���y���j&<<
0$���4[G�D�W��^��DF    IDAT���צRr�f]����^��]8wF�4Sߺ���r0u�$�H9	��5�pH�&�a$�\��D��0�W�Xo�l�h���u蠘٣����7lz~I���
J)͎��}R?8+С��"	;��u�(!kF��P��l?������hH�����~C=�˫����CJ��hC0rr�z�zd�=�t����e[[]�n��Z2���t�h���*��I�*Q��p�NY��)�<24l׮�U�!��x�����)zl'`Gd���\�!�9����"��8G�1���t�BgҚV�u6I��S�¨1�3��W	;$�#'�3�]�P��yA����8����%vU�}}�YO��ZH$V)UZjO�k��; �����g����{_G$�U�rqadh�z������@���Q/rb��VV�;�#��-�M i�T4qZG1E���d(��%���T�� �	#���4f2��P=V%;E	\+�S(����(r���z����-���6%N%3kH%8|̫��9H/�2�q����#������������Q���U�yȳ�Ǵ�?�wn^�&!E��4�����s�>�ۭ��M�Y3���oNės�viM�E�Lo��z��t���|Th�@0$�H�f����2���z��&���v�� u}^��@��H�":
�:
���F�跑��78��0��cdfCӊ���jk�˞f��S8=5j����r֖�����
<�K��{'G�U����o��?�N��μ�\wk-�l�����&�����*�����-�zu\%=��dA-��D�O�l�Ha�	%-�� �=�������� 	7�e�����@��^ 3
#�L�S����!z��ϧ�N�ق��Z�}�[��c�����Y|I܌w\��m���1$B}�����`�&X�������S^���ӧ����@���i���ۿ4�p���7;0$Z�4�ԧ�y��E�=)�K2�|��%ϐ�ږ�ˑ�qŌ ���J `��Q y�E4�:U�u��)128$س��؍7���]�c�
���>��"4�R5��S
��G`������:��*�\w��4�O����PV���l�i?��ٹ3�e��=�o��T�s������4����M}c�8��	����DHE�H� I��[e%2U�%K�J�R(YU]6�-�TI�h�e��?�*A� A"q��;;;y��g�s�}sr����wW ���5սݷ��}o8�9�y�s*�K2��D����?��B�ᵚ>��i���B�d ��.��D��<H�h\,�˴��/����[v��{��gG�m�]H ��?�����r�Ӓ������;��ւ��ոM�@��I	ԖXi�_)�c��&h5�����c'�=}o/@Rnym�ff�T�Dӳ�JXK4���H��҂x������%���NY�ձ��9���9�r���~�~H�/}�K�ꫯ��S�{PO���C����I�H����,z�-<�S�����+SbuuUk��2�:<M-���c�l��,9׫���6`(Ѥ�x$*{�r�
G��IT���D�s	S�<Pǵ�rH�ZN���x ���g#B�_�%��/�g����3��ݛ�}��߽q{�/�"I�Z*5���DrŜ7ٱ0���Q�!�J6�|�H6���%�ɤ�K:���jL#y�qr+<f�+jI ����}׻�|�ŗ^�͝m�|dK1��̤0��U A>y�
��mi"�'��ja���J�:M����������>�����x\�x��M�|�U���AS�;o�OyQ���/��WqK%	�U�?{	O�����������|�bS��2�ja���o<ش�7����F��̨� �� �(�m�$�E�5�̈́-�A��%&/��H!G��)�|Ҝ$�&���ڴ���]J�ae���lfy�B�tZ�:L�Y�$�;;7-�j{{�^��$ɃV�k�6e�������]����h山�����<��J���"��ZQ�<i8c��o&�¼���������@r#��WA<�ژ���A�$�M7��_�ꎏ�2ܔ��$�:��/�R�?8:�F�m�ts��E��#��j$U�p��H��@i_���� �z/~�l��X&� ]Xأ�a$,//l,//�g�gg�ׇ߯�����|+ߓ��}��_�u�����_oE=q�(����\�Hͺ�G)7N�1n'˚�$y_@������i���9�xDG=a�z?���M���A�����z����>g�6��W��;v��}ߧ��%Bn��%�qO�3�P0����T��|�_x���A�S��y�}|lm����~�c���|B����׬�g���qRȉ�^C����(��%����6Ꮤ��l�5����E�� �q*�+�D��m�m���]�y�v��e ��U�������7��E=��OMmԻ���� �����,f#�[.y}3�����WU��֦���QԀq���lzi��fǸ���&~,}kvv�D���ŗ_с��@�2�aV�j&��;���a"l��>�k����KJ� ���u^b�e�nR-T�� u�Im2��Zx�懁��؋Rߌ�{ָV�O�b 9P�h���'�$���ef�z۳�P�qt|b'О�&
���h)\�u�%T��˫�t>y�I�
&A�7൨*�u��-6؁sg������ե��X���wS���V���{_�ܬ޽w�?|�ʵ���;��D��(�JxWN�2�"W�����dR&H�]&���)R��c�D+N\�P�0���.0a!\�kw�
������{�{�����M�>��ڋ:��
;���$09Ɔ��a�A�{��N_��$����8� �'4�6��+���?�{ꉋ�q�g^�~���5�]a��/��� ���Ƣ\��8b\� r老r����fE�!����|�&�xU��`�'*��ѱ�[�o��lg��N�`�H	���+�(,�"#�9�<�	��?=�c�"�h�����1)�(O��̴0ȕ�U�Y��2FR�'yH<H���=��ڶF+����e��T������(d̎�lok[���kj���K���{\ڬ��8H>�	�	ZB�U:�]��<<H���|h�p���������,��!k���/��b1f���K&��o���Ag %�&��"-2�)s�9Z\�O��ɤ���m��RRL$Z���Tf���j�9.=��aJes6̒��k�6�%��h<��vjfg�6���}��;m?8��
�S�ZZ(a#r��fmiy���s�~�#�������mye{�v�ƍ��z�����?,��"�.�_r�Y��]�PBV+0�p�o�&��O��n�= ]+5�
�><��0� ��F��Hi�O��^�,�L�f���Ab iz������?z�p-j��}x�!Ҧ����qiU��M��]̎t2BC�Nv܋2u:
������t�-�h�l��C��'�������z�%���7y��sԏ�R�Ƌ*`�%�Ҽ��0�%�����R�	3f[{vg��=|�e���� K��f��A�&����S�.�1)�L �.'�`��`�p�>3xv�u�<vV��v	x�S��Tw�ww�v|t`{�;�&�kai^���0<��0���}��ف7'p���/}�������scFI!b2��-2�H��a��x�Ph��T��g�8�Ax�a"�.�h<�u3<H����8��|l�a�7��1Ȍ�*�/���)��
*���r�F���u�6��n֕�_\^�A&g�ʴ�U�J6T%�鍻0�cX-�/��I���|�{/�\j����M���Bv����(qeq���v��c?�������^�m �b_�s翼q��_=<�b2���������z��!%���]��9+TK�y@�PR�N*.��i�]�����r�%��P��a �X����� �9y>k�j���w�S��ύ;��� �����|�cS�������Ϣ���l�ͭ��2�0����%��7W����~��Z�;�{�$���w-'՜�d�D�I8��'Ec��2��`ع��Q��J�W�}2Y�}$��z,$%�D�1	9ܾ�n�6����i�NG�����R�̍��@FE�Q:�{6M���,��<J��9�3�"ɼ�9��-�b�U�J��8���	���vH����Ë��r��hB�|A%���5HQ�~l��V)�������~�N����`���B(0�TJ�Ux�*e]]����ݭm{����N�ʶ�rv\��8Ɠ߅G�{8�ei
��dWু߆!�$�D����Pu>�kj����ã}]�����g���>C6��j�ݦ5v��:�A�M�Z"*�ʴ���8=//r8ʍ3�|<z���bð{���o�ś�+������	�"!��a>D�mqa�֖�liy��s���쇞{��3��kז^�y��=����G�LH�&#����l =c�a�d?�	35��x�%J
坵=�B������� b���&�*c�jz� r�\f$I�[�|J���~�7���;J���`:�$����Db�������=����@�1J'5�����d�#���w��Ο[�nwdw���/�dZ4�����L��� a3�	�1�p\,�rY5�^�^Tx���m�6#�:l�:��H.%��:2f�v���{��i��{�H�\%XR�2ӽY؝��Ȃ���/<ǐ|�R�F���[X\��\\�:fF�
R��Tf\Q?<���mK%j�V��ck63?+�N�o�'�͓#H��T��n>�������#S%kuH�6Ӂ�w�θ�ֽ�m]Ϭ��@����_ZZ���%yU<?����1b�Fv;�Yd�����CZx`��g��}B�z2D�=��c�9l�g�9��7�.j\�|%15�MŰg�Y�qh';6�B��$>Z�ZevѲ�Y�) ������L���mD؄ؿ@2ac&��P������QbGJN�]Yƃ��������sϽ�=5�/޸�?<����|� ����%u�����0y�Α��P������1x@y��M��%:$]��^d�*�	|��>�T�X������K
�̆bړ��x�q��3����H��q��iL�@
�S�m�JY[�"�+�,�kl�X�Z�ّ�%�S��qOpD9K�8c�����{�kϯY�=���n�K��"U��%�	�&��k�3'>7�<� �,Bƌn��iS�͢�sT���ڌ͖�2��SB��J@�bL/�m�ڭ;�%pp|Ғ�$��u��j�ТvY^Q�i^T�#c�a<��x%�h��¨������U�S677+>��ڪM/̩~�X�Y�d�Ž�q\�ݝ"�f�̊J�
%��5�]!7C0�H]��#��o~��H\ 9\:�"ǋ���*��M�<{��?��v��kv��-�yuզJ+�]x|<22�ѫ&�C��a������=�x��z���b��0s�..���W��yD"��7�a��u����ͺ5�v�S?�� E#��	��h��̊5�(n(�ēV&�:X�À�� ����)㎁$�H��#���=	%��P}F0�ڢԙ>sf��_������z�4��v�M%͵{�������do��1d��Tc���U�g *���SJt�T��6�Ζ�ǈ<V��T��v�'�T&�,�[$�8GT��
���NOK�ҥ't�_������#�r��	����s���BLI������<[��L�	�&D�.����P��*��C�1�O>~�Z����׮�@v�}�W]�x��O�4���"\B.�g�:�LU�R?G���a����cIĸ�+���h��pk{l ��ͱ�89A����g��9WXꦒ0WɃv����F���#��nf�V9Ge�̌��Jְy�����t	I�M8	��Ⱥl�<�S��ݪ[�~d�Q�{����o}�2d}a/y���>��ApU<�C?$1�?�#?�
 ���ekw�6=3'6�%�C�K���Y��"��5���e�o6���Sr+�6�F(�%+��Ai�j����9dt��ߞ����}klY�h7�r��p}�K*��Ι���~}�b3s�V�8������k���PC��a��;�O���΀�x�I����¯>vv�/��w��6��7�ݷ�?w��)������}��wwv�g�H��1丄!��D�F�wګZXa��햻�)@���@�[+�s"aB�X^�����Bo�T�3_�Ե���%U���g��S��_�@� ԏ�x*��T���I�P�?I\C�$Q�[&�M�x%��7|���%�V�۵�Ѓ|�)�����2��U 1Uq�X�Xpl�����c�?,̎K.�C�G�%���P��驒��EH�!�|wh�`s�$�c`��fÍ5�#!��JwR�,!p�5�i<݈v%-��ь)Ԁ�PKP#;ҁ2�� ���d��sVN��T�����><���-#Q$��Vln~^,����1���uZu+�3�A�~�w���'��	�����IR<"9�s�:A�#?�v����� ��s�l���ZÍd|"�/�����r9EP��0�V�(�*n$�0�al0$!���unG�-������F�!вa�ĎwZ�~h�ů�,�<�\�A�&9,�� [������^����&Y-�I*KRf8Ly�b���^��KI�!�"r}���@2��\V	�3K+�����kg��y���e�m����|����x��w��S��T�m>�!B����W8�d�^�!��EfJ�qr��H'}��f��Fx\���In��c���aG��JФ��	5ipE�=�ve�է>%O!�DfQ����,�|��ᛥ�9I=
�V��&Z�� :��#�C�[�*I0�U?�w��+|�;����W^�~%���>�����Z���Hm0I!Ce(�P'�n
�}��8E[�_ԽD��7��m�y��=�"I�Px��0T$�E�Rm)P�BB^	�:��EW�籰5��>*a ��r*9?/�r~q���d@2��ww�D������+6;7�u4 E%X�V�H=��m�����ٵ7,�$��Pu�ɋzW���<QI��G��?bxx�ٹ�AݾwW�l/�j�Ć�ψ��#�T�+H<Xv�06��Rio8Zk	#/�u�q�x�~����%T%�b��}���VӺ�{v��i�֡F}+��V#|R(�lT��ly�F�iȑtG����vCL�S:�m�D�㾵�R����\�u��k�u��*e���c�,R%���,�ٵ3�����W�g����(������������褱�b�Cۏ1ᚺ��U&�&O��`o=�k�(~6�;*�@)a�K�.al�T��$�N����Bޤ��`b4!��#q='�%+��TQQD+��|�S��[�o[A|;����b8x�M����s���*
�ݛL���Y�U�8ߓju�+L�­��hU�Y�ߺf��ݕ�	�!1����Rk<Ê�^�?�H66��,҂��!؛���Ey���Q�+�!��0fv��}�u��O��h���zu��='!C5!	e.Kv�	�!����w\�K�Ϊ�Jw�Xm��I�A�����*E%kƥ�T���n���!����H6<��j�2�x�:�:	pO�)��X-��`CSG�Э��m��D�I:^ؙ�/@�)#6�J?����H�
��G��j�!>��XwD��<��T��/�pB�/�]>�y�nb?�b-�̈H�aQ?9������$)#4��r�Y��Ȏ�6�xo�
ֳ�k%�I���3�/ϚM�ذX����T�$�
�J���z���S���	<5��ddJd/t5�!xJ���v�S�3�03MC�����/+�zvv���VM�m{���g_��S���O��{o9>9�*b ��Zԉ�^����t�҆�M*N*�Qc��
oI��Iwl`$-��g��    IDATW����AQ��j�1R���ث�C�o�Z[bά�IՇ�]�_�f�nOƅg��G	e4J)L$����3�6�6^�꧊d K�4�B�=�/ϕ���AR�!�~뺽~�(�LyO���V�s;���.g��F�Ja=�'�ϻ�yN�k)?e -@ҿ��Q��-�6%i8| ���#�~��Hԇ'uH�R�M��6y
�b�A�3���K���c�a��ۮ�^=Y�ϙN�!W�US$ږ�V��'R ٢��ݶ��C�z�)Y�V�fcr�$��6�~�͜`(thK��/�	i�[�N�]+�+��Һk{�����ǟ��{�n߾�N� ^|�Q{0���N����?֖���+�dŸۣ�\�X�����]����u��p�/�{L��=>�~�Zq��Y�Ty}��ڶu�g���ur`���F����<	Z�N[�P��T�r�Y��P�����|y\"��d�Da��dz�B&�5����dH-�N'�rG��Ðo���O/-���?�?��ojG��]������[OQʧ���hޕtڠ�p�(��s!�HV����H��t���ˣK`e�GN{�w�$S��r��~xj��N�Z�!k�ĭ^�B�	yx��Y�L��@���V/_�l���$��a|�H��cd���*z�8B���OR0�����z=-Ha���H!ȑ����O>e�x�;���xDI��Ƈ��s �f`|�T,ja��#�]��0��9a���fJ���g�ӶP���b1��񰇼�ȣ��ݼ{OU!Ɠfӎ�F �:����!wCI��$V5&a<'�&��苬�B�TZ��Iz)�H��u�	U��S)��������}H��q����@*���x8К"yE�l���~��"%%i���l�������Fbi�d0�癧����˯�ZM��ʫ�ڣ�h�����RS���5�i�sx�l~�W��?�3<Q�,�.72� [ad���_ҡ
���-�,�Κj��cl���8ܷ�Mt�V��[��$��嚍�S�)�Y�:o�ڼe���JN���DKJ���#�$_�N���Wu]김�֚Z�
S	6?W����wl������rq��/��O����3�ߑ�|����^�v�o���n��T��$ǜ����0��A�����e~|��Mi.��b���:Pr��MH�����W&T���s����Ł7
�K��1�XX���Q��j�E(�����N�u"��%��(�__)����AF�1�T��DIX�h�E�S5�T�� ���|al Ϭ�I���'.e{V<�޲�1!C��J�^W/Jbbw��v��Z��/Hz�,�/J�P�;b�A���}dv��ʃ�K�e��2�$�: Z}����8�&qrؤ���I��0�����#B�����.)��AE��C�j��h(����w�A������,���ă�s/U�d�N�u�Ɠ���ݲ[��hY�'Ͷ�Jx�u�@�J�]�n���}�}���-�W����CNH�~箼GpIheQb�q��V&��9��cKu���1�����$?�N��(	e�Fu���7�{{;�/��N�32�Rm��y|l��}k�wm4��t�l��3$HhNU�m���@��+�ʕA�8������i��I�q2b{�)�ȁ�� �њJ�,eR�xy�`��V�N��K�k�{���̯=��S�g>�3������w�~�޿�yo�}�f]�x3�<�sx04K�fL�U�V��:��j�Ĥ�~{`���l�N}�xxT��P7��3QE8a�� CV�obNء�^�+岭��H�g{o׮���ݽ{o�A���O�2<Ye	S��AF�>#�b��s(�B��7!v�D��I[Ҟv;6?;g�|���ɧ��t��;��ν�vD�.D}KEaE����@�'7uJ��gg�Y،�B|6'����	����y�<i������֝�je*u�V�`` Y�
�'��4^:8��ԉ�Jz��kK�X���=�kO��Fz���F}gh�I�y}]m&�R�[+)���d
m�`�+���[w���%�R���F�^:!1<Q~O�LFX�|��^|ѹ��K�Zk�Ymd����(�y�͝����'\<��:)pG?@|��u���}^�|�yG����c2�8&ڈV�]J���6����u(.hY�sl���D�d%t&�8�l�ʬu2Ef+��8�I�x�\����]��F���1���v��T��h#]��e�1�9[Y��j>k�NÆ�6�����̯^x�ɿ���|��w�@~���'o޻�/nܾ�� �J`0\�s�O���E��R��A���l�[o��� -�$f�������Fe�6٪\NxS�v���G`j<I�0���Dm���)0H�N�nݾ#�Hǩ���^ϫ0 z�4]_1�
<�I�N�4$E�h:Q#����)S�07o�~�;�ɧ�Ե �I�6�6 ��C
�H`�e<�}1�R�S[K"�̠k������W�ux` O)�~��	��ݺmw=H�t��$Ć��s�����0j��0�bj�'h�#ÞJq'U�=PH�t�凁��#]1G��xm>z$|�����դ��OUR��������O�Ѓ�����?:-���'��C�Z���Ї� ź>kfzNM�0�_�r�5����a����˥��A�%J���@2^��c�����#l7�l
9*�*�0��}��w����z
K!��[�7���Y�=�)%m858��X���k6Ȗ�G9f�h�W�%�?�B�{��X'G�󟢏o�A� �F?���%�� �9[E׳���k�����V�����k?�џqr�^�Q����ƹ[����k�o�(�j`u��C�AQO��4�FYEzK'~�։�1&$�4�R�aQ����1�tNx]��g�Ó��Q�!&���Mm7;��a�1z���rȊ]�~C�Q$i�6�o�@�%<�"ʪR�$����У]���u���qCM�!�b�dl6��b �x�	y�{��2���#�wg
I����]�ړiM��=�ʫD��(�� 'т1Mu�H2�+sj�2���#���#��~�<��8�AF�-E�4�Ȑ>c\
�T�v�qs�Fٱ=�Y�Tr����{
�	��:�qI7�8R����jM5��sV��N���Ӻ��z��{�8���#;>���)�..�!�O�eR��Y�t?��?h��[��d
�I���Í*1$Y�b�w��RZ��U%�(�u�x��〃�^c`��gj������<�S*�e ˥��xW�6I�!�K��l�mZ�~`�Nˬ߱>I�
���vd�b�����6ȕ-W����S��
[L�5��K��P�ЁIG�=i '=H%}�N[N�3K��tR���A�sӶP+�����i��k��p�]\=��>��O�|��;�k7����W^�򓀽T$�}M2R�_��M�B���S!Lg���j��0���g���9"�5*̦�3�V�A�~W$s�(9�דj�#���ua���Y��=����>q!_z�=�կ�y��WI@m��Q�h����:0���kI���<ɔ�o9h��l�ww��y�۞�K/Z�Zy��-��ߵ�Ɖ0�)�J
R��� �K^�6H"�GOj��4A�%;�I����<� ����0��6�l}s�vw���i�I�i��cO�h�y�&j�yΨ��i�
�PI�7HQ�� ���U������s�$p����7��d~G�
Gǚ Z6 u�^GTW�<)�ag��\���_5�.��7�1ƣ����<�Μ�ٷ>k��+�"j������Ϻ=�ϡ��~z���xW���#��r7�b#�aKXnHa�z���}47Ɩ<�*�"N���z��	��m���a�z�c��u$��oX&O��YefVE�ڜ�g-[��Nj�j�\��~�0�Q]*����̈́��O�f�>��多V�!�dZ�9�I�Ns�ڽ��
�mس�Z�V槭�8����:��������ǿ��H��[��̃�ys���w~�ڭ[�{�d(T�Am�|Ҡ�L�����C��C��ŀj���CF�QF���Ne�
�)����
E�h��0�L��Y���LXL�<�d���^vW��r�Ҁ��y��W��y� �e ���nGx���k"���y���Ǖ8n�y&Z���~�)S���'�g�}v��_p�6�v�Z�o���sLț����~�p`�d$����р��PB��6�$�,ұ(���Voh�7������	���P�q�Bp�vI|=�I"i�N�<�6�(�e��ͳ��9��,q$ȥ���gt��Ab��Yo5�0v���.��-�����8���pA��7�ʓͪ`����=�D�dOs�|C0I��[N���]�ؙ�v�-�mme�~�Q�(�=*��Dƕ:v ���#$k��ϊ
4���O�"q z�{*�"$���:#8�0U��;.G��<iyo��в�۶Od {�Cy��ō��/��2%e���Sz���,_����#J[�V�Mk���"�,,�S]Ȁ�"����3��׳�F��yA��_�	�CMo*��j�`s�h��EK �{�O=��_�������}���wd �<{�����������J(:�P�B�^�qJ�HzeY���vpt�J%��.6�����-(ɨ��2��Tm��Q�-#�������˳�����#n
!�;��.�׮\�{7�h9�Ë�v'�Q� �ǩ>�s���Dҍ�K�Q�%W7�p`cAO���49�����,σ�>z��M���'��U?���Gym*���!Ov����S6�|���	�0�G�Z.�T7��۽��hY�׵�����hޥ�O���,��hʤ�B¡X7fkC'�U%OR���D�S��$�1�D�a	��{���e����|$��W..(:�Ѕ�¼����&�C��f�:�I笗�9-ȓ�T��A[�%u(z� לۧ?�i[�_R�WX	��Ç���x�$�ꕕ3kN#Jk�q �
�c�~(��$��{��S!�ā������a�  Q)����H���v�j�����;6ja ��>2�$s���,W"{�����03U�Lq�:ü�5�0���f�1W�M�W8i u{��pF���W���{��?c�+z��V+S6S)�lm���wd ����'�z�/����=���F��f~N�a�+_��v������� k�hud ��.Z$�0HH��){���8����B|u��P��.�pJE�+��~�j-�j�E0N�����wxv�g2�IN���Xc�Yп�ߧS��.�˯��LdT�$O�:a��E����{J?z��u��
���B3���x��H���`�o{����!����k����=�ḼN�C�.��&>G�#��[����Ԣ�d Y��=;�<�uؾX�d�}Z��x`�Y����ݽ}����� �Ɓ��A�*cBS&m��~�q����H�� 4�8j����Φ(��+*a�g��s�xYI���]��F���Ж��#��;��|>�d�~�:QvU6)�N�7���=�_��eϝ}L��ڗ�����{��.�x�q\���hjx��d�Ȩ��G6������"����s��S7�TpDS���~0�1�K<���E�z�m{����^+d G���{v�s�sCdV�V�P�Y/S�Q�l�BU�cn�j]�J��:�>���s�NbmD�0�b<�j>�|�p�YyJ�My���+��L�b�5*�
�vU9�lqa��s���������=1�\��Ç�[�����^{�}'�*�o�+��33�(;X���U��hZ�.x'N���Y��1߁�����Ԕ��'mdHU��w��b�b�����#	D��BA����}�'��׮ڗ���ڄb �R ����z�`�8�I�&ɋgaaL�����@�y7�����``d�/�� .$X%^����=���W>��"�8A.K�/�FA�w%^��P�3!����qD�linA�1����f���6w��Ɲ�:!Uom��@��6�G^s+�'�|-R7Lq�<�-b'2��q`0��;�jp�Qޗ���������>�ە���bΙ;�N$��c.9������tJ;%3h�OTG� :��3�O{�-�U�����M�cϟ;�H�^4�?z��}�j���k;��63�=r�#�3�����_Fm��C�j�8�e|RYgD6�oߠ�~P�Dy�x��H�����f`o���=>��Y��Aܴ<�k�6� �Y+�PR8m=*����6ʖ,_�Z2H�'�W4�DE��g/�:yHjћ.�b����ĝW�9ך�*���Tֲ���mR�0z�҅9���_��?��{f �Zoݿ�_�җ��Ύ����d8RS-�c�&���$��x~M��f�,s�4H�2�G}�I�D�Cj�	��p�>]}�{����Ғ�	A��B�
��ps˞������v�K�a���A���'�?j�=�.����6�:
"���{�mgϜ�f�>����B�������g�Q��.og�kfԇ;rJ����@ �XT������Ԭ�+vQ�mGU ],�ʵ�Vo��1��HI|0�X�ҁ���Qt�$2Lb���1t�!.��R�A����+ ^l�D���ֹ\��<H0H�t����Ɨ� y�QOv������?���ζ�:܋��i[
oc������e�XH�h�R	fLm>�n^����x<rU���x�(������	�яđ$�֝"�� �(�Ǒu��8�<���{�{�"�z��"��e>�o���6_-[����;v��i�v�rY�}2�ˏ��:�h�9*Fʵ;�I�l�rO��m��Z���|�Dpb}8>�˨'1e%v&�\��c��,�%>M��u�I-�����4rب{b��]+�2�g�}���VV�������Y�o���;;gomo���_�ڿ���C+��Ur��d ���5�������4�!&wlВ�-����6Tѥ�%�:5�E���D}����fS	���A7A#NB�I�L�W�fo�p^a<���\��-V���V<�!��B=%�X|qB���/�����{3����y
�yҰ��bΟ�7Ǐg���S"	C��eX(�&��h��\N-6|��x�Rk�Zᒁǐ,�{�
8X媚&c�������ׯ����5�)�`�{Ca��0B������g�����i�%���;I�5�X�}%�.�� ЖJ%x��Ϫ(�<���`Ŕ��Ƈ�-p��ޮ*��'���'���N_��ߑH ��������4�+<��(��9���I��{E�bIq$�b~�b額F$ͳ��B 9�G��a 'a$d�2<(�'<�ςX��0I�?���g������N�v�u�c��m�z
��勞����ί*k=��e;�����^vۘ��y^��f���8���S��`0�p:��
Aq��v�.���a��^�_(<|�?����e�}�6���p�z�w��ٿ�S���d2�V�M��;6�W���66���+����1�S��x��N<�a^��	���!��xqx�݁g�Cl��V�����L�@d�z�S���坦�P����ʃL��t�sj%Jsk��id�:��Z  }���0�1κ�+F���l�(C�^_�M�Nmd��Z�.�?[��wArl�k��F�g�`Wf�c�͔�d����B[����]�@���)t,�u��>!�K҆���d%E2�3�+W���[w�R��ѐ�oHZ��A�\�)��<H���$�N�� ��$!�b��HS.ci�4��@Vg��%�.2�qZA5QO 7pT6��)hg'�N�H$t����1�����ă��r��[�i��������.���9HNQ��g^�qta����;�3�h/��bR�$G`���G�D������)(��@
kO5��`���3T�Tb43%��F\d����=>�n�к�#��d�H�em���]������    IDAT̚��������� ;%��L�?Z��J������:$��R�d��$�-���=㫞�ݮ�C�� �L�PjP^����`�o[}KY�J������'?���w�K��k.�z�࿻z�Ɵ���A��ZmF������IspOB_�	a u�I��=ʷX��2ZC��g0,�a7��n��F�R%9�I���4ô��{��50�L��s��깳vcC�H~/�%���K��&D�\$��� ��h(��YE��z^d�~�}dh�C@7�k�I(Uxy��l���6Q\�����Fo0���:�u��@F�
/�g�3�K[��Ug�0��s��mM2ԯ]�n�E�?��\FYl�a�es�^Ru���Կ%<��x�R/.�j����B�Z�I��("������!��l7O��z��Hu�d��/�{�<ؐ�N$�81���;�-O�nz��s�)5�E/ x�Oj��	��\-W����y[�_p���k��g3�I��R�=;;m;;{�ۿ�y�r���Y�H��x-�>/W�KJ�_��0�Q{-7n̡�7*�1{E�%��9 �]����Fr���e�Ɖ�������9c�jѦ��.]��̒qX�Ȃp����)~"�B���O�$R�9�^J��n��#�M��q�,�6+�,���9�����������k5la���Ͼ��?����or��߱����7sc���������oݮ��(V�fHVس�x\�.�dX^�B�Z�sPy.��|� �ᩌ���槐Ts��K�L� �m:�I�!3B�&eϐX+�X(ip	}�\i���A���x����;��v ?��9��fMm����2���I���a�����z��j5����T�,�w��/\|�h#j���BI�z���FCO0 y��P#�v���$�R�i~�U6���Q���B��甬Q��.�����ݽ�nۻ{� U����hh�g���)��h��^��ٓ��	锰���qݤX���[���ǥN���W�w��zMu�#��
9sK&��H���s����M��9<<&n7������ho�^�D��mi3G��	,[t�^ߩGsZ��3�WF�7���ptx,q�R�l�r�v�w���/	��uG�W��)X/�ʡ_)<%㰁��u�J��6Y�unff�leyM��;_��5UFضѠk�^��CH��u��݄�Y�v���E+��<�Ӓ�c�(ݡ�5D|}�d�-��R%�[����LI92�c���	��OAA�̈́�@T���i���AqL�Gsv~�"�j[v�?����G��������*>a%�s97�_�s�ۻ��7�*���<RF}���C�Nx��C�v�L���A� ��<Z�D�0�2�+U=�l4lV��ry�}��1���$�>n�h%ЊT��nX�u^4��.�k?�����~���¥��/��[n�[S2`ORx�0�!?V����T����q6p#	�J� ��J$�6ciy���=�X,*̂Bx��>��)b|��r���/�R�:���t�`3����/���7�J+�������T�#k �E9�ҩ��TT�������Pc��$yG�<Ƥ|�0�u�gq��(իo.��a k�Xj���pc������s��tHI����j*��-;I�d�t������^|��<�|Ɩ��� ]R�ω�@�A��$V����c��@��{�Rj!�xpx���u�5T�0�/\��X	CyJ�'��8g��u�g�S�wu����%�/~�kV?>�A�#��hбr	�rh��&)�>�+�V�K��&���P�M�_��+R������so�&\�a�aK�_�}��83-�4ړ$�6�5���=����U�ؒThI� �Eh#k�f]��Jy�����_����~���.������}��~���l{s���r��9�_��GƲ�vj@?�.�30E���1��i��6��%��<p�Ds�SAX��ffPb�w|��m�˂�6��q
�����J�#ܧ�飞<D�{V�y�x鈯��=���ڋ�/��;w��+�$�NNN�K*��n-���tJ��,h��$d�=m���7p��l��wBi�IB�͇!Գ�ę�)d���$<Ye�U'K�w*Ť��>���L��n�CXV�!
TҤٴ|&c�V׮߸a7n�R�5�6��� ��FÐ�`��	Z>I���+/'�Ë�W$o¨�I:��T�*x�U����J42j�y �ăý1^I���r2&����5u��ݶ�z^�-1�%v*�a>�;���vC�M�yZp%!�1klvv�Οw�X��DՓd�8��v$��D��#�&�ܺ-�0��m)�����A1D2�(��PT�NJv����2�{�}�͠5�T�)� �Jvq��!���"#_(Ymf����V(�GFp�c�0M!�ޭX]���USvƳ�9����.�!^�<&JZ�=FU��o/*�p�^O$أ��� �׽dt<�f���NP$�.����s�-�����O��^F�b ?{�ڇ���ǯ_�������~< �q�z��J#�G�s~�P�5@Z	�ě*+�,��(p����Fh6�cn�ctJl[CJB%k")��OEh���+4��0�!8���>�ڏ}������=��KJ:�u4K� ��i���K�� ��'�M4��@�Ru�K��Glt�N\���άx�ʵ5i�NOۥ�/�J
|9z�DR�E����KU`��
�Me�UB�Z���6W�J�dS���;����W^�͝$d�N�	"�A��&rRB���J����؊�}�%or�F�k�T���O�E*?f�=�Q�td�V7��It��;�����0���,��u����ߕ�
k��*�Ø��{�F���P��̿0FO�y�$ggϞӜ�+�,��8�-g̚7�\�H`��}v̳�R�X� &č�#3�#%?SeW���D%S`��gl�o�K�C}th�!F>�]��9��E�#�1U����z�8��7t/��$z��	����$���)�'�)��{��&��*:���ƀ�{&bA���%	�n���t�t����_~l��_�Ї>���ol&�+�7��q���_z���V�GQ�T�k.zӰ��4)��AR��F�,�iF,W�0�)0̶�t�wq)��n(d��;���P[�/�O�%TS�V,1��F)"5��{��K�C?�!%F��;���ξ�`�,
�y�0��Z	Ӧ��a�$H�B�D����X3�x�(��8�]\�W�˽�6��sgTK�Ǆ�]@�c�� �o%���T��!�����@Q��ڌ2�t5$�&�q,9c�6��׾��ݸsGp~ƦH=;�� M�Q�y�y�K#�y��
�P_�-n�'���'�9��A��UL���1�M�3yaI6�챗����)q
���r�<;'��+{��S��	#�ѝ��B���z�<?��7{)�u�t�0�G���R�R��ǮC�E1�io�$Zq�
���S?���RH�5�L��If��p:	�#Ϡ�2hd��9Ur��w�5��.M���q�&F�<�,���!��:��΅R�k�b �^�Dz����m��RT%� *��
o��!�<�)�H�$H�S�s��!8����`��ү{������s���'>�S_W��ͦ�b _��\�}��߾r���׽Q<�<�5�����:rqO�Z�{+9��t:CQ�Y%�؞lv��f����*�`H��JI�4iBR@%tZ`�$�0T�����aF-���Y����=j����ו�h��2���)�2Q��*��ov����
M��:����N��S�*a� 	6�H�+�2��*5B�լ
C*�ӼQ�A�M�Cg��=;��DyƢ�0*����fk�2��|�P��ؙ�(nm��/���8���$��"�%�`0G#����Y�ƃ�I�\5��"�0a #t��Q�88�ޥ��Z*dS��:$�ZO�F#L6�1O��}��zO<�o�8��OBq�)ZVJ"��O2v��H�b�BA����Ӻ;{V:�Q���(1w�%��Ί�#�&�~���U�ٻpt:"�2=E\C��	�N��~�����}�V�d���\8���JF���JE�4�v��rP������ ���CB���X��1l){M�3E��G,�Hv;e�&�x��A��~�R��wl:ᙨ,�}Yߝ�F�j�⍳�K����o$N�=1���ʯ��g_{���{p\���������a�
(����\5|֓Q��]ޢ��W�x(��&-ǲ���Y�c�R;������^,�B�����K]	|�!��$�oZ��K����m�p��ܾ��-��l�aዩ��+Dx�'�4#����%�y0d�؈\��q_�yf9���8$�Ǹ6��%�|R�B���/�[���Bڝ�S�d���� 좋�{��J���M1C�4oQ�|sln���˗�ֽu; 4$��)��b��yv�~�ݶg#��������𨃩4��������F�R��P��/�6��k����3�ᕒ�����3J�5��wrt,B��%�x ��0@p��!"gO ��> �-V�%r�̣�s��%�UK�$8�H���Í��cvL�=d0Y0�7�i?�g�o�*CG��8��c43?D܋XJϕ^c������[����k����Y)�S0�mu�+i�G}��H��7��Eg(�ړ�f1�rT{Z��x�t<u���ļ�A�����y��u�Q�\�B|o=R��2�۠svu�_�9���~�C���o6����o�g��|��ݼ�K{GǫH^1��c%�Xsz��6#,���}�Gz�*(��&�ũ8N�p��ioa�v�D�#oச]���1q�Mxs�r�^��&0��`��TYA'#�}��t߻�6>��i,\�ҩ�K���R[��Gq=��f���� �yh�G>[�z���}�A�9�ll�͝M���e,�XF5y�lD<s��,>�!Z��ϋ���kQN)dA+����܂�7EQ<J�����﫩���5����J.xN����޾����YFǧ�&z���߽q���3��k�ʰ+�B�Q,���d���$X��T��3�~j�)2��z��hj�B�&�wj�ަ��� ~�� tOΐ�ﵻ�'Ɓ�axl��̘��# ���7�&�$�y<����IŜy��k(�K�DX|̜��g�Eɬ$P�� ��*��T�$i:pO�=JZ��+����F��V�F&/x�J %�8�R�cT�@풧I�>��h�@^A,R��6	!��RJ��@P�N����8�7�Zy�1��n�P�X'���Ν�O��O����Q��{}��o^�����[���d���UFu�5 P	��ޠ�`��Z�R���V�%��w*��zC V ��L��.h��Hϋ��P�I��FN�Ë,�/ڀc�j2ɼ��$L������_����Hrl�r��!GR�!�ʠ/`��Ԥ��ֳ	g�ȁ��\�>*^b!Ȁ�0)��|��������vii���i�.t�����-��W.�A��/�d�h@�P� �)We у,������_����Y�\4�$$&u�N�^j"�w �ae���3���.�IA<5W#���p�H��&�K�U�9��MO���K��qp�=�yΒ�r�r0�ǇG)�L<Qh-$PRͷڄ���yr���'{�T�"ƏC�p����P-G����������B �ԞX\� u'�=}��KvU�%.�n�4ǎ���ҩ�o�<j��(@��h��oυ�I��H��*;>p�/���u#}O�F�2ρs=%dR6Z��y�s��;A��!IT;�	V�&��߯fM5�?��=7��E) yբO�p-0�j�C�Y-���٥���'?��o(L�=� �p��/��¯X��������y��2M�\�������E�6�B��7��c�&�}1A4'RmwG����P<|K������h N�k�u�^6�7U�i�>W��RM�r�*��� w{mi|�9�j�~������=�x�Y�)�G�8/��0�,J8l,2B0��I�5)�8���b�bA���T�70^8��52����p��9� :�9� 
r��w@۳�#�IKͰ8�f��q�Mol$��r �C�����.��uB<'�bCC�/H�2z�J������m�F�(/6~�<Ȥ,=W�� �q���\��8G�]d�v�2�89Zښxֵ��+�6� $2���L�&��+[Ͷw[��:�P$�z>���p�y�S�ψ���/i���'�y����{飌9QB"�G�D(Ѓ��`x�Cֺ�)"�ԱP�I�&R.::�j�\n\��0�܋�Gu7�Rm$�3�]�z�.����R���-��>���:CfN��Ҹ\#�)�UBǩ{��2W�����<ǂq��d8�`��@5�崄�377�$eu���l��W��O�����b_��w^~�oZ�����{���}�E�)�l�~�����h���'��d*�(,	�Z$���X㎓MSQ���5�2��G�>���k´ש%�	�DR����qC=F��U�Z���<S��j���t8LΞ�}�����:V��RO_�{RHK����e�q�`�G��I��̹kR('���l���:׏�ë��I�/1�2�M�G^R�W�Ab�O{+�F�n�3��ky�C�!�gg����-�4��J'3�u��}��l��e�E�\�{�����*�^<�Hz�N{���8�qSH��Q�z��~�Z�^�O��A,g,���M�#;�Vqye�!�9�C�I��	����U��{�Pc
��7#ʠn�d�h~�=t�+�g>Y�:{K�84����o ���
�'��ԜN	$��VK*�G�c�Q���oP,A;��jNi-t�MU������@�a��:��;NT��rN�rז0�o�RA�Q��3���8k�Wx�j�R��R��i�;�%z�qZ�Av/TIthkU[^^�ZZ^��3������~�����z�c��bs�O}�K8l��Ǎ��~����w-HqV�Z�k5���&Li+�a�GCp?�TE봽�2^�c^��/�S��!�YA
o�䡭��H��r(6FmEDآ����4��΀W�_��Ñ�#p.��Y+�������<5v��E�p�6�T�'�d@u�Q0��A�Qu��C�������Z�$�B��2��3���E�C�F���Sx�ͪ��9^;�f�Yd�����[iÀ��հ)����0gkK+2�y*���IT�^���/]~Y��i;ۧ�E;��)�ٸ���@j�$#)��$y��$6&n[Z��w̱`��`���� �AO|�1��@�r�<�L�'�NY��D����l�t�tP��۸�ȣPaaaI�j�ю�����eQWR,����]�;<������ �)^p�$��~�֣g{�� Ð����Qg�x�ŵy� <F�PI$����o<E�e�Y�t��z�+�*�aT���0��g���JX��b%m8px_�����`0�D<��/��U����'��L{^b�r!�tC��_���;�<;I��t��������տ�g>��o(����@�����7�7���o^��wﯟ�AP�`����e��kڠ�i)067eݎY�<o���q��oO<(@j��Լ��OP���t�j�?~Q�
QU����<'1�����@I��[Z������i1��bU�,���'��O?#��r�5�eCV �u4�J����F�_R���wJ���s:�s�Jx�cxR�032�x'd�14x��ƳԎ3��e�Y�k$\/��Q�&�ͩ�"���F�"�@�P�v��]ɣ����PZ膝�:�;�dK���ؗz�$�	�kx\�ôS/�]+�I������q&���c�'!:졐́�DB���f=�$Bн�$��C���l�T{6��̷Z�VH�8�����ʡf�%��2Fa D~/�.�R���s��*	7��դ�tv�'6e�S��G��#�����+�dW��<�429<a!P����`<8�	Ԙ�B�*�<�yV�!B-�3"`}0��%��Q�К���z*�l    IDAT D;C��'��\��]��eR��\i7t�-��3,d�|�>�a,�^WޮC��5pM'��!)q���`qq������Zy�_��?����wՃ���/\��W��7��~퇦J��ܨ_�:��z��3]+�sVE���5o��:�\�j�|��C���r���X�ԂBG�#���� -@ҿv�/�Et�n�M�k9��� 3�x�R0'i��Z8<8��æ���X3����,v�p)JH�mo����}�7e4C�@�4��m�h,
6)��{_q��"v��o���\xY$*t����c.�I���	���a�r�����#���n��EO�� r��P��W�}��n�)��~|�:lpX�.�_��6�Gv?�ִ�G&+��[ �WEJO�%�cy��L.#�9���ҡ�F2�#�$�\�F>'Ulƅl5*=̛B��͵�����H�膝�-���u���Ҵ f�<��03gO\�d�\�"H]�s�='5+p)`<X?a #�uM��S9��<&&%�|}�
�����P}6�M��db)��?��{羨��pI���X!k6;W�Ko9c3�e���(��A�=��P��H� �FW��оB͉��f�k�>ъ%J��R�0F���a���*����5��@U�'�D��X�Mjj�wm���n�9{旟z������������uɕ����W�߸{�#�����tufЫ?�m^:9�>�����s[^B��l�Lɺ팽v��봒�-�`����NI\|0���VՃwui��>vF�_Qa�s�����۠�,�,�����@t��GxT߷HŽ��Y;�kڃ�[v|ԶQᴰIM\�j�.=n�>�v��W��.5p&�WlD&���B����T�u2p���!���1�����и!eA,/;N��;����D�q������^�+I�p[�3Y�4K�sJB ��­� S�Ckҽ�#5���%�n��9��:��Jt�ی��ԍjx���ŧ;U��BF�6̆��� R{X��[)�����^}v����0���L%o���v�g�{<��2:e�vB1��m�����'�R=���E;:���ܬ"Z�ZG	!ad��)'�f(1�5?M,)c�ڞ�v�CL5��j�p\
1�;W�$�}	��kBao:�����1$Q$@Vc<7S���y����UQ�FE+����w��kI�5?$�ڝ�������݆�P�b�����7�����K�����#f"ϑ������H3�m�u�ZJ�œb��Q,�n�OOnme���+�����ֿ����ȴٳ_�v�Z�����������������D�la���<?�f���}�/�Çvt�ڍ�ُBJ�
Y��\^Y���m��襇Lϐ�C�)�f�������Ў�����߲z�HR��B�fg��޵�Wn۝�T��\�u�~�扖���P�c��í�2v�XO����
W��)8ayFN��	o7��ʸ&��ӄ�{4,���9�p���9��85%��Ik�	�'Q���AXg����U�T�_Y��Xl�&2q'u;<���//�#{�ʌD����IX���8��-��Q��#O4%)&�C�Py���pu��A��8b��gf�4]�}x���Gh�g���$�'�(��8�@����B�͸�R&+�q�Z���՗/+�aFd�z`��cny��4�ΐ��+�{�8�16*z|�{N��P{"�J�����K�����!pT���(y2�D�L���_@�aa�=� 3]���%{˹e+�r6]�RY.�c��]���2]$�=xp|�峖�Re�NN�s`;�G��u`��'֢=�(o�)�`����Zj˽��D3�#��4������*�)[}zf���j��6U��6��l}������o�{f �|��7�m���{�����Z˖�(D��M�+��٧��o��Q��z�!�.H8H����~Φ��j�IwyqI
7�<'�s#�NK����Jb������-�lw灍��U8�v��6-���[�Zm�n�|h7nl��ƮM��O*�>��Q��ș���3o{V�q�`������0l,4�I��{XN7���������P*L`<F�J�5Q~J:�Y�$��QW�<����ֳR7�:"��ؤjʋ�h��+*��Wjԝ��ޯ�|��V���:�uŜ�q�y�Ix�D�jx���IB*�����ǵ���O�g�{���+�@� ��zy*c��8]��GEW$NɢdP�Fĳ����DW&�RI��뾿0�T���{%#��Qn=���	�����0�~�J��ɍ�:�I�u�rE�X���J�e�X�
u3`�)��;��ϗu8��!�S��q�Qijߓ��SXX��j9ok���<k�(fe�҆DSqiqN Z�B��ڌdNy����C�`TP2�j{u��a������o��vU��|guJ<Iֆ'�Ph"d�N��V*�l@�`�m'��-���s�칿?����K�ֿ�o�H�;3��Ѩ��y����_�o_x�螄$�']{��M{�k�Y&K/�i�_X�riڨ��u�5��s�R�t�')jUZ]q������
jfq��O��>���G6к�p�a�����6:+��:�b;{-{�yl6vm���nnz�O�*AU[;�jo�;�!�Ee�g�]�lܢ6��	ۊM#� !O�= ����r���	g{i�7;�BΓ��{�v�\2�i��c�ߪc��f��6�'!!s��y�~���cJL�i=�ݗ.dvW1wq���E���&�HF�5@��*�k��戰1JNc�����#��J��BN-2�7�$h�Ȓ���6���Rm7�қ�O9�I��h���P��y���+�O����x���]Dg>�_�1[�?�#���H����}\����u�z���<�Yt�(C�a0��ma�jsse[Y��Z��%��e�=�������M^�J��)1���� �;�r✲�E�����N��_m��=ą����Q�,�]!�L�VS	g&� K�
ՙ��'��ߞx���>��k߬��f����@rCۭ�?����ם��W^{�6l���=|��T���\�3g.Yuz^X��� D��q>g�[�����jr�b�c��C�ڕ������
�4<�͇�mEP��C���vToX�3����9���dl�����ٰF�#OVa��|�T���[�j����?{�dk~]���~�����1�<�hd	c�!	c���,c��PĔ!.��P!�]�P�B(1F� X`I������Kiƣѝ�;�νw��}ީ���u��)lJ��Ҫ���>��|��_���^{m$i:�c U�*-o�5S��8e� �J)�U\]��2��r�j�_�U�Es��jD@�z�qȠ�\����*`Q^���$��b�S4 �O3�HNN�q@�k�)�}�`���/Z�J�R�F�����ϯ~��\�� ��u����$W�
5�cR��D8J�5�"A�/w��(�W����"@�'�J����ӗ��)�I�m��W�#��T"T76_cg�o���cԹ�0��E�%sh�g�5�h��zm���`{�� /�ad��	~��#T���������'�r���v�¹�1�d�&;���T h@d�G���������2�Ѥ���;p_��t��u��mۭ;��{g?��0�_�E�G��C�AM4�3��)eD����^�e���|�{��M�B�����������l�f?��g?���~�#q��_Ѵ�v��ɫ�K�����{�Z��\���_�E/�3p/��<�*���t�Q��t�\�v]c&���8������9ܿW.?{wn*�"��u����N&1]r���i��j׮ފ���W.?#���%o�+�q�����k�L6iH^,jV��LѪ��w+ �*o���\Y���ecnv�Sp/����F��q���p%��C��)v�4�� $���*wI�S&J��|��qj �t=���*�0��Ա��O���QS$f��j�e���R+������{S�X��SF��ylLY��M�T���s���8�eV;�0?SW;^��f3Z�f]��P�v�'@S�x��������������xIm��x��>s���s;�wAF��ϟ�o�%a�^�ˠ�����~+�������]F[�U�?.�lCedߴDȀU��*�-�B�=�z3��K��n4���x<9�P�+�[���E?:��݃�z�Z�x���uy��b�Kd�an+���x�ν���=\x���雾)-�>�_/(@�\�ͽ?�˟���?���qxp+����o��8w���7c��Il��}(�z�	y �w�=q���V�?�d5��Z��n�؋zΤ��8��ٍ)z��7�еsK�k\cv�ISi��f%&�UQ	�ŝ�����W���������m��7~]#I`��r��DW��v�֞/FvJ�s��:~���^��JT�E��s����).<~�,*Gg�粘�ECx+��2&��KvmTA�jT
Q�\R,U�O��դ���d�T�Y�td昋��Rœ�zp���V�b��HGۊ���e8Y"�YUۊ1Cf�}���
$UDO�V�b-�r�X�t�h��)�d�K��k6�*���8���a@��:�s�!N�닾�("����M�� ��t�|X��.x>����S��T��u�0�x���E�یsg�e0{p��N�F���Wz��4 )�t��=/6jߣ��PT8��<i��ֹh5S�FԨawe�3�t��2��:���T�y�����g����)�܈A��__4۽�[[;�;x�����Mߑ �ǯ /^����?�+�{��'�f�щ��q���Ltsk'�3�$a`��X&��x�����O=Ǵ>q!�8:ޏ�0�����X.HS;�޵��)�HK����e�M�\���/�����Zqpx���Ph�E�]�ҥ˪:��U���b���{_�Ξϙ���9���P��x=�oHE0���`�~�i�:�� Aw�<�E��[�y�:�S�%�Q�����1t�~,pyP��g�)�R�E�(Ҷ�7w
r�Ѡ�4 ]_��-�)�;�~�N熋_,=�J_K����=/��j^��)�B
� ��ˉm���;�& ����<�y�Iw	�[�2%�!q}"��<D�D�>��.��J;��� �yU��(UgΉ�++��ޮ�"�j�MZk��T�LT,�6��j�|$E��۸�gW���3Z�:6�����!bsL�R�Q����+ޯݡ���Hk�����)ĐJכtqAiELfKu��G��d�Y�
 �v���)sm��gĹ��-3�����?�� ��ưm�b�ys����˿��|g��/(@^�u��/^�{������{bgk=$L][0�dA�#)��uck�z�+㞻��"�����^�܎`V/ŋ��vF��yVQ-x��<�w�.�h�j��T�ԥG�e̖���K�~2�'����{����<h��������bx2���8Ν������� �,�0�.�>IHEJm3��CL5��s9=2��k�p}��"�*[�� #�+���n��I���B�� �r��0((�toO�"ڦ��Ru���8��bR.h?���ҝ�l�w�R/)��JD�]s� y-Gf�S��i}阑�e����b&�R}�ЭA�W�)T���������{C�-��`&,�p�Ni�l>.��I�0y3%0UA�#F��U���f�N��Q��_�j��a����$���qoom(ͱ��w���D��]Ω��Ǥ����9�U �W�G�C'Eу�ц�:@�V�Z/:=f��b�@�����hP�-'���>���Xb���;kR�Լ�G�7�nY�P����W�s�{\�'iY�ȵ9��̙�s���w���1p\��
�����r����[o?w�l4��!a(��O&�P���{�ɋq��F��:�899���;�`�9>8؍�,�v-&��Mi;܉{�O'���W��t3\g��������T��1Yv��"RJ�j�b>ǝ��L�ڵg5��9��#?;Z!�Y���$��߳�{ɔ55i�$/Q��~ܤDl��ܬ<Ǒ�ݺ"^����r�J��d�Q�2���rn�c'oT@����X8�l#[!���g�o�PI���Iw�6.�:��5Կl�s�(����j{��$O}
̅� �e�!���^cSgk�p�[�Z��	����i]f��9;�4�=�I�f�4�k_Ml��\�nO�շ\� �b�H�Bm+	8Fs�������,5]��`�-�-<��摠�Al�>���!;�_�|�=�H9�y܉��oǃ��?6�#�3��q�L�� $��Œ�3����J���d_-�:�zW
���Z�WA�@3b��-�'�kW �i����? �cP�z���HէQa��7��)�;7oސ��i���t^�5~rs��w���z�7<@^�ti����y�����u��5������C���ǝ���{%�G�x|��)���=�f��LR��;�w�7��AI������?�X��o�u��-& \����1�\�z��9�Jڍ��|����
 ���"����Bz���<0SK3�1���z���N4���K��(;2B0�A�8x/ �G����{�ޓH����<v�(��[K�����jl;6G�Dɹ!F��,��M�s:�qj��V
�i#M��ү�苒�;�2˹A̮��e4�|��9�9^�$#�<?p�FdED��R�6��B��;��$��w2���k�G���R�2�r]�*s��%���)�V��J��s���� �9�Ƹ�0k9k�F	_oo�	��'�<���p�	����+�w��w�����E��Lw�l[[������8>�H��b�ف������z�����E���F7�N2�e�f�N'�19ً��@J%�F��AL�u��肚4jщ�\Ƞ�s��f<��\������;��7~�����_��S������R�V�����,n�~6n�8K/:H�N����lE�}�$� Nw��ZJ<��7���J�ř��_�~%�^{Z3�Y�3�l��֝�8؛�d֌�3�E�3�TD�-N���l����ĥ�����;PE	i6�����lT�i?D�Ǘ�8d(ܘ�J�L9���kv���M�H,�qTYM��oϻ�#Qz��㿩\W���u5?uxx�(���>�.��79�A�~�?�%D K�x1������e]�#�lE�j>���ŧ�)�#<^�iqFhXni
����zÀ+u��fc�����:"�b��g)|5�/f�q���j�2��*C [�d���2��U���u37i���>�-�.I��O��2�):m_��F�f��k_"e��|&���/w� ���A|۷�-���o��S������	�?R��tzw�@2+�Hzr�(��#�q��}1��ɬ.E5��Ƈ�H�i�<��t/�'�ܓى �YQڀ[��������k'K�{^�����z�{�����^��,2|��^��c��?��F+�z��|�&�iz ��;�]�8vKq�v�ܗ���zZ0!�˘O�F?�l�љ�cnU����ݻ��K��N>�7܎��R���[�Q�6v���T�p2U�=���U\{�F<��GQ��p>�Ϝ�O�Z����K�FV;�dG��k���T!HGj���� �5J�>w{���"�ϑ
��+r���%YtiJ�s`��@-��~29�󅞰L�T�p��5sh��"a�95W�}� �� j�a��l�3�~p�$�� �E�^_�S_H2�_ӣ h�X�4S]������1s�I
s��w�T�i�N�ɗ�]5=�x����1d�s��r[�ũ �WnlY�������]mq��&(��kx�A�#,s�{��B'�������{�Z�7����#��Xl�{�����gj����VLN����c����n�U`k4˽pt��qt;����(���Yk;e�tb<>��V4Z���V�͹4P/95"~��i��?�蓟g\|q8H��ӟ����w߳���n4��p�7}��.e)�ǯ    IDAT���/w�������Y1�xx�Ǉw�7:�>gH�J3� S8��N��i64����ٻ$�y'e�up&�!h
V�+13m���N��ޏ��_�����cv�j��\$ R�P��"�N7e7D�J��iv+0��تv��<sS"�=�~�X��v����#��I�:pJ��B-8}��?��q\v��F(^���on�b ��x���d�	���g�U�X��pt��A���,�\�8[W�K��G��׬ȑd�""���(�\nP�\�fӹqp �AW�����*#G]����p����)�/zEoP~-s���O�1���0ّ�S��"�>��U���IK%�#̒h��!Eƌ�5���y��C���x�����{��mq��V\|ⱸ~��\tp2�i�rP�z�����h�W#�	W��,�Q�c��	.;�h��� :��P.�b~��@��d�d��)���Vt�C�{�͘�^H?I��)�b�V��Ho��}��]��A�_��<��t�R���|��}W��#,�n3(Hv�L�;R4@A�x���A�U��8:ؗ�K��KR�L�֎/��V���2�۱�s^����T� �q������
�{�@B%�칻b9��>���O?ۘȞ;�90}��!���Z�n+���F�@����H���[�h`t�]]�<���ԋ��o|KJ�c]�a!V9-/>G�Na��
�e#�^�}�@��2���U�*�&1I����S���6��J%�\�8��ռ/_�SY�y��6'*N�K[6�ż�ע�j:U{)<�Sp�{����)���i�"m�e*F������K�Ǧf��>V��ӡk|vo�byw�(}��G��<*��7�u�_6���N���PQ�ۢ��sN�\x���8쳉Qܚ�d	��^������I�'7�_�;�o�~~T3��D�V_
 I��a�����F?�ntc�ڳyS���" Y��zL�����c>9PT:���s'��:cviGLޱY q�b3�F�v���V���������������$��S���릋�{"V�c��6J͈^��[}I
H��ܺ)���yr�	��p ,�'9�il�[F�Vu9h��0�\pif��ol�pc+qi9�w{�3q|4���\M�Uov����qr<��s�_y�bl�=gv�E���!����D#�6�����]�[j��	�x�REV�)��� �Z��ׂ.��^�>Ud1�(����c�!?9b�u�Sl�Y��I��ez=Q��[ꐽ�c9�F��ˋX�J2��hO硌�t�[��T�Y�px Dчs���96I�g:>��3�����td���L'���Lq�LG��<�xS �o�<�* 7���^�V;%�@��=��.`*��ρ�MF�Tn��yX�#w���>w )�F�m��  9nsج	�ܙ!d+���r�N'G�~Y����-�^!��T ���w�ߣ0�B1�@,��jF����t����?܉���f�X�:L9�$b~�v-�}��;���b����lZ�G�<���&����Y�����p���}�����}@�?��o_ܜM��>99�����y���Qt{����f'q�w[d��!Q#���2&�̴A~�����2�a6��*f��>[\���t;�F�7vo���d:�aoX���蘾�nt�#q��x�ҵ��'?#�3g��hcSr  R�,\HfݔH�x�Q�֙m��H����:J?7�i��<�7O�
s��� �(CY�P-8�r]N��D�(J�AW�ǝ,�8�'E�g�B�Oɼ���oU��}�I- C��)��9��Px*aZќ�S�Bs���0>���p�i��u�rs�J�۽݇�YYx?�DOt�p�T�$eUJ�N�B^[�R3М��-F�:n�׋��ϐ@X�K��h՛���tQΜ1���6�%H&0Zi`�����E������\؊��گ�������7����j���`%��ҘL9�h�G+�&3���N3��mBQ���yp$7-�4�u�XjѦ�����m�u�_1$V�ޔG���� ���E������{����������`_/Jɧy��寺�{�o��xr'�F[��!mG�i�O �"�^���Iܼ~-nߺ��4�SҠt(�ώc5�m�p��@V�q�ވ��ާv�X=M���}���	�'TΎ��w�.=�T�܅��3�I�[�TK�A�=ʔ:�e H���,����h#7�=�L�@݂����{
�H�H�<��*P��*����aʙn�N�	C�R��I�2I�4@ʪj��ZGY8U
Z�QdO��P�[���rj�ɢ�g������bʨ���mM���'*�3x�0ӫ�0y-' ����8RP�]��*���e�-}윇u�WRP������;�uG��\���Jʎ�gpV�_L�HG�~O]O9���Ǝ��."e ��������&�+���[��__��_��y1��PU�y3v��s����dG��`dA�;���Y�SZ	06��@0��3��m\70�'��(ĺ�F�)0ѣ=&����P���埶�)���:�������������h ye���O<�ݷv���zc�A���?}��б���dq��n 8ͮ�\04q�E6�X��==��s��1��֊�ƙ��>�V_) }��TeY$����i\y�ٸ�의L�Y�ۻ"��Μ�G%<��K2�O���#�ں�q����d�~2"#��(�dN��ڲ�V���qu�P(*#̝��T�&�aF$g܀\��"K���Y% kJPi��k�:��F(���RHl� ��=��r����)� �$�)��9����V�#�&Z5��y��2GL��y��A�%޺�Pg��u�����ˠ*=ŋEq�)t��#S�^Ց��˼�����75����-�VT��.��&��$����P
���$ݝ���߻��<��}��+_.;�.�M�&��I����M�̞|#g�c�C��l��q��èՙ>���K�~�����=X������c�Ym��@���!^�Z3m���{}�޺���~`4�o����G)�Z��EH�>�oy����ڲ>yM�E�%�,ZMҭ�Z�� ٟ�|E$;��4�/�haº���N����w�����f�ϙhu7��H� 0�j�=z2W�荛����O��k��6�>0�^ds{G�#7*3�������.RLݨ���t����%j%��n��V��&�gK�ߑ�3@:2r�₂��
4DD ��A�N�"��h.����|T 弸jC�W�Bɕ-4���pQp�7�_7#�,`X���c��K��p�σ�MO�����j��$%Jȼx��β��~?:c�iP��]S_�~��#�o�f����gA~��ͼ&��s��d���p���i`���z1��M8y���4�\͊�X�c �q��hi��&G��;sf3��B�ݔ>��Mt�����h��_�v2&j�h�F�鎣���:9Bp��c�`�Hz����8~U��s�"uιXB�4�9���m�	��h�R�?z�;����θ���b�q/*@>|���?��_8>��z�ΘP�D����=ۛc����ٍ��zJ�#��?�]7�6d�u����y�j�fSU��E��S�nv��ۈVg�F'j�~�V5��i=����ãi\�~3>���bw�8��q�mi$;�A�#U�u�;9R339	��#nqs]ڧ�)�F��7"��&����|WI��ju���Q� ���r�<���5q��bJ�l*@ɼ!�S���HifĎ@y�QB���rZZ�`�(�*�Tʹ��1�<����ܜ$Ȥ�|os��YR�J#�S�����y^]���c�i+��|���
��%��
}�M�Q�M�4-��Q�c���{�����T/8?*�-3������h|]�,Du̳��ff����"�j����f\8F�G��}("��� ��wU+  M	�QT���1��^{��M��s:_U��=t�3f�3P�5.?D������"�f�c3 )p2���h�v����㷾�[����_�s^T��`?���kW/��f+����J��>i
R�N����l�[�ֺ����F�`�޹���.�?�$?����(���wc���3���%r�P������bȼ�g,��rV��zD�V
{H*��.l�ˍ���$7O�?,E��ֆ�'RVb��)WS+��+D��iUP쨪EV�*")Wc���
	�*Uo��@����>���ge�w�N�J�@��A�9QW�>K�`��l���C���Y�����������B�?w�vK��r�t��~��#Yo�B-T�2Un�	��F�g���JU[�j鐒|��"����Ϗ_W�ǅG��B5ŏ�qz��tO��e<nc��N��<O�Y��?T�Z�dq �ߍ��-Q&T������P$	HB��"�\A��)��.3�&���;����N�� $E�T) �!:�v�����`�ظތ��Ta*��$h�C�z�_u���/P�����E������'�|��L���l�b;5V�&mH��K�C���S����{La�
�j��D���W-�<ژ�C�#�L��x�V;ڭ�Z�]�O=�tܼuG;�}v-+vM�^Fڻ�aS�b"�K1�V�Jy�W��|t��i�
`qQ���נ�JVM��	�J��*�%:�o $�_N����iVh%� ��O�!���tǜ�x�z��LcћZ��Bw�����u9
tԽ��ӌ���|�|^�n]Q.�)�"�{�u�K'	���  ���%��9ȕ*�)pe1�`��8�ѿ�������l����8DG�V8���9���JGv�JL��X��k	�T�8��*����U��2�,� 0���]��k�� ����i7e^��9R��35Fn�g���*�L&G��8��&��Ezk�6�� �zӯ��sV��ݓJ�Y��:G*-N���J�(2k��p�q0��x�x�����w}�L�||{����G~��׮^��e�ߘ�8��z�"܉��V�����Q�:�[����|�1ȶ�c*��M�5�].9�e���g��X��k�8<��͛�q驧Uucw��k����."�ۮ�9ϒpp��
�4��.m��"m�,�Ĥ�2Z�S�*��W�9,/Ҽ�O;e\ ��H9E�W$(J�KŔ�N���32a!�o��tܘ	�m[� ��ٙ�po?n޸���Rʅ̤���;��&92�>-���l�1G�Tӿ�41�:��E)b�m�X���6�Q=ǎV=��Հm�te ��� 5������A��8+X��g���`�Z̚�V�*_�"�7I$��� ��B�5_��6�rO!�I�5�� �	@,7!�ۦ�a6��Nl�p���xԏ��@�;6K4�������՘K���%s�KE������N��D��ykBs�;�����ْ!���.{�XI��=ĉ G��G�lm�����^��@�� �'�<��ȧ?�gw�X�W��^[UK��!1p��(���p�~`D�k�7bj�n5���q����H3��
H��i���Gγw��-�5y޼��e*�xk;F�qt��h����t<W6U4)��ѝ,2G^8��M^�Dr-/c\��s���@5��F��&Y(U9�k�S��R�Uq�,��R�#�Թ���ͱ"n.D��"�����5ۛ(�x���Y�J�R�E�����f�7 ���]C�l�p�Q��JG{Y�(�F֙2k]���هWR^Gg#ܾ�X�J������f�� m��l~O����������r H]�z��ju�Jd�cHD,3vʹ�:��&����- �����%��I){���CO5h�[���}��fln��&�'J�� �\.�rÊN�� �T�]3F�굕I1~�h��i=���X����b
%��ߑ�uڽ����?�������o}��Q���@���?���{����b�!.ۓ�p׎�RNn��7oޖc�UKۤXE[��"��sS�I�XM�v��0-X�Ƹ������߼}'��.���lD���y):mZ벪iW��Tou������6r�2��Ǌ@/f�b��<(J�2�=:���4HZ�����.~^<]��&�E�7���fd��� 3z@ ���r�6���������pG�GZ�s��4�k����������l�6d�?W�_ug�LPIa�"�f��`d��z�iq
թ���m[��̓��c��-�������<;��|1�MwA����R�S����s�_��Ѡo��lǛ
�6�A����]c�k H��*����~��[7S�Iۚ�����4E�}�W$9�w4�~�Is �@8�����TlU�P�p�׊��;q�v���dD�5����6b��v��?c�8�S�d4|rck��}ə/��/�k��`_2 ��Gw~���=���^���h7bs���,Ji�t�hA�\��8>�-$#�>���0�~w��3�'q�6�bw�8v�c��8�8D�6#��>]4�톽�7ӕG|a�����tm�˲�DGʹ�"�N�(���4i�39�7m��fW�1�#��~��r*�.�n�F��9,�� ��4j}�`x\q�_"�Fv����� �8�@�MT�"��94��N�|�$��u,�G�Z��q�<����7:���W>o����u}�Y^F5��\�J�BP�+��u9f�[1��U	���������Z���q�l��y@|�M=�V8-~��\Z��	xs�o����|�z ��Cy�|ߴy_9��FT�j�2�8<���#OZK=��2]�Ũռ^�s�ۢ�ƛ#q��^W��t/��#�#��ۿ��7q�	 �l�,�>��j���#b[m��T�nun�9�w�;g��Co�ƫ_�h�W{�@rp�����3��ר-��䀞ሖ���Ⱥ�)����V�8ܽ%�8�|nxE-�44m�GE+�y�Z\|�Jܸy[��^]�}�ifuG"VnƬ��X�A��2�g���?�lvu!jP�LS�^Z�\�H�����|SW�-�'��p�����Ec��s�yS/:G`�T���g���F����$����sD���GV�i��Y��� b�����Ϸ�C@�4�UMW��������o RQ[I-���&
.�sE�P��
}>��"�U��p��j2��1v��e��(2�)���Etfy��Wf%�!f�JW��V�K)��&�u����=� uJ�{%�6���&3�H�U��]ft�0~��NS���:yM��D�x�1��x��/Q4)�qQ��4F�n��dA�-9w̱澀c�(�L�I蘉��	��N�X�5����C�;��������ਵ�b����{��ŋ���ʿ�/�vo���ѻ�Q��|�� �� �
�Z���Oa����pO�1�,��FG^�r5���'<d��T�gs�F���͎E�.�ʥVz��,���x�bf��T�Q����T����xj蚧���G�N�v�����>[��B0G��f)iU�g�� �E�\x<���=��-ڬ��΢ݣ����uzɴǜ�)fz.j��z���v�J�YS���D���xO�>��E�v��X�Z�:7���9Ҿv�&���Hj2�-s��8�vnD��k $`�MS���3��gO�,^<߼��h�9b��`�|s��T<��t�u��F�w��:Ů�T�\N��$h���y�'
h����^�$�R��hP�����D�tN����q�]�5�W�n�\��Ad@N�q#�)����@w���x�z�*2�������7�����+���?x���X��HN�����y੧��_��[.�s��QT{�m�ư����4�o���-�U5�1�dO=}%n��J~0R�e3��xF%�xR_���Z;�8�L1L�k'/��%?{֌#RlER��f�r� I�E�'/^���G{�;
�B4��T��ҭS�2���<�*dA�Z��\�=�p�A
ܝ�eOn:��|p~0d�:�K�h�]�P��='�Os��''�"�R��{Ǔ    IDAT�؅�|.��R��C�O]�'�Y������A���>�P1`X����"�(cjB��S�r��5�I�[��J���']+�I 9W​l)�떑��O�p��*A���6w�ىSH^���l�{=��7Y�;� -E�oH���CMЖKD�Y��fUě�wJzD�y������ƨ?��`�^;����м��E��&Y3�ن !@޿f��bՊ����J&�7���V���ό�������Ͼ���� 9���>�z�g��}�o�����s׫6�R7ȗ��� D��?>8�k�>W�\Q� �$����>�V7�4!bڃ�鑦��t����t�8�r�B�Ud���9o¥�����5�E4�㣇ܑ���j��S%],w���E���^�-J��U��NC���3 #��DIa����ad��/����h�998U��E��\����ˈ4��C�4�VӠi@�s���{G�.t@�@k��}����T�32���Ħs��[jq��ae�A<�(�Ϳ��q(���{'��%��ŗ���N	���J��Jn^ќ��ǀ�i�����ڨ�	���% �%������T�Ag��)��6��g ڸKq���|��X�W�O���Y���B�g����3�i5��li�Mz�c���B<]6{��~w��~��=���=�PJ@^���\�9��O���.?��_G�wk�̖�z��e�*3b��|����d�ȕ�Ϩ����P7����r ��BKW:?W)i(]+Bgs8 �o�u����� H��2���Ӧ���+* T ���c�t��:�5�����������s�a�f��;�wF�%U+�Eއ�рD����yq(���/�s��M1A/�N.X8uG����|G&�8};btD�s�M������ҳ���u\�C0�@�2G�G��ud�".���eF����&�����5�&�a9�5-��Vf"����`_w���	R��f] ��U� ��)��s��;���O#fm�eS���8��xM��%*����5VK����.P��t�$��ފ�Ο�s;8��t���Ѷ��xt�x�}���uic8��F��#���jg��ܗ$@r���������loo}5����2ZB���G?�H��Ň`on�`c�A\ ʑT){��7�s)�@nP@>o�SwJ��`p\��r\���$�����"�2h��Qmre9����O��K*kq�#sm�����]�/ ���;<X� �H�T���Gá�?G�U����9��It5-���� �&j� �c��E�|g�<� E���vķ��@��p��N�hCq�ܝx�8��h�ό|L��L�%@ �͜�{�r��3@r�Y7
h�.̦��#L��T#I/F�îE�����71�#����)�7mr�R`�=��ӛ��M*ɊR7+�0g̘ѻ��2��M,��{�":�u��������M�%�"d7���_��2)���$�1��l����}Qdl%��o5�?�����=]����/Y�|����/^���N�]��[�8=CO����+W�ƕ��'	@�ʇqs�����/E�����&Btq/�o��3�=p�\q�&�K�q�Y�z���%(ABsc�"�L���M�Ss�$�%U��W,~�����F^0,J��z~1��^M����2�7�Vͦ	�����7G�'h�,=�Fr���B �Y�כ*��SD�}��ZW���ſ�5E��
��́�����-��3a����R+d�+ >�?ȯV}<$ql���E+�����J�q)rT= Q4��S�%i3��ޜo�O]������VYI?9���S�e���E�������,�N���Vʀ�m��Y?�����ࡴ�J3E�I�qn�9�-�Nt�	�����x���4����M'cX�	��H���xe?�l�H��.��x{�m�d9���i��V�������|��/fj�s��H����+��k��on7�[,Z���'��'�|2�ܼ���,<=���9{>��}w���ؾp.���A�#+�hKT���~'_���)Oq��ѓ�-��������8�S
.��P_�>el�Ac2Ϫ"��u%�8\�U�Kin��UԺ�gJ$� �D�k@o6���L(�*>�v��pu�B�zh���4ۂ��"�nw�U�QJeP�[>ZzM��y�����J=|�Si�)ǩl�����V��(��=\���dA��%E�\��@FsP*�G����_u4�nzd*Lx��;�D	��'�Q+u�I"�9�1�S&qҲ��4�����	vl���c�r�}��W�|n���&�����qK��>�T;8�f�S..@��)��_�D,^�u'�� ���wrt���4\�~�N��U�8�j>�� ��^���ڣ�z����-��-)�x��^� ����/�^�����O|ōk�nܼ~��䵧�~:n\���&j�X.����w����n��=�%�Ӵ2�MCۛ�i�0и�H���N����A�i�#���#�8P
JH����Rvr��H�Wvh�����:k~q��{EE��,�*g��xK��`�ő���N6G���VF���U�j�C.�\�i��� 2��Mǀ�ݠ�� c����%r��j��<�{cd":C��J i
��pDb>����N!����X�]�:�~{S�&��ip�a�Rk�FIx�VG�T��.{Hu�hP�TO�f���	�˵��� J��bT��ֱ�G�������I�*���
O��/�[咨�� 	��<dZ=�t\sl����/(��P 9$��K�j6�O7����{��~����=��Ar�{�c�K�?��KO=��;�n�_�/�>>�Օ˗��^�ǻ�j�#�#zo���^v_�Ϟ�\G��f-�X�KK��nƠ7@r��U=�o�5^
�|)����ԋ/n�鋒��
�(U 5��ke,*��#-`n��#� �2o�"\�Kq�P���Ε��~k`+�9r��킈��ۨ� j}��� ��u�Jv����U Zα#1~v+��C�
��|'�0^��]4��KY�'��4F�x;�Hu���%��"�]�j�(�S%��7��S~���]^�|O=���:�(�-^O���,dXb���4�DSw�@[6���i��s*W�2[sb4]2�Ko�PA��f�5`�=|%u���b�,�e�U��Kv��.��;*<\Pծ��g�::܏)�PުȇRAѕ!
 9��o����>���w�?��w�+�֗��K:���\�_��/�=���OǏ>���Cz���V��_��2̬�=;����z���;Q�bȉ^1oBdtA���Ƒ@�ŧ\\T��|C����d�kh����ˍ��su^�y)��뫤lH��9�n��-������7�u��'<��o0�Xx}RlGj�<��?]���T�{n�:m�uu��:�?�,�)�SX��j*���HG���:ٖ��KOV��@0Z
�����:מ��>���f�r�/���07K3�����S��tT��N����N.�8d�k�F��g�����o������3Cq�J��xޟ\�*@��ܡ��>��O�n|�z��K�Ʃ�f����6U�$���Q-���]���i��w�V�ɋ��Y��4k����Q_>��x��x�ǝ�x�;���2����o���|��/{泏���o>�����?���g�ĠݗVK�,��X��G�}����ڊ�$�h�hp�f+�d���wLE�L�,L N���捷��ý"�I��b)�ͅq��"C"�R����reҋPN9��[U���e8�e0*�5���x=�ږt�HR5���鏢��)�y�����g��*�g�t�Tޭ�4�U�-�S�VƤ�'"��Qiw��*�9N��7s<��S�<��7�l-���� ���?7�Swrof.ܘbP����H�|�7��un��w�F�?-���#ZGi��&��<Q�ǝF�P���ozk7�����
��FՑ�
��7Ҁo^S	�2��3�^a�B:1[Dm1�cLcnߌ�	��1�ʟ�pE���7Ʊ��}y�����l�������g-��B=�7@^y�ѝ'����=�ɏ������v����`��EN؍W��a[܌z�����;��0:Tg�X��Wc<��e��"�<��L�ޖF����
�o���;�U�8�?��V>)�(E�C�KJX��������vwn�2�F=�t6����ѻ�a�� 	���s���ZM�%�7��@�����Ź�o|vW�u��c�*Mr���-]�M
��y�b\�>�b
�>��=��L�MqL�����Sqs�,����3���wͧ��f����'�2����Q�耢o��3<�,j�;<ZW�l����n�Hs���
�kP��%ס��j�S1�w��Ua��VZ�oE�Y:�Ly�������~}�Jω"k���ڹ�w<������7"��F���~��Q;6�9�wzt���?>�>s��n���+����_���?���� O=��?�����g>�W�����ot&؟MO�MI��zO�ZXc�8�<g�ƹ{��x��q,��hQ-f�t�H��]6�\$A��´I��w}sCHS���|k$NK2���+wy�ڥ9�R}�1]��y#D�Hxn�N�<�:@W}-�eU�C�"����c�� Y�N��Q��2p1����ڎ�>N��azq;Ք{t����4�iZ�?���W�C���y�Y�qa�E��X�r�Ș�	�*VmN�<�#��M��[���6�}�Flfp��\l2E�&$0*��U��:�(������|�PAZslJ�K��Q�ߛ'@��SJw�Y�\�c8���r]䵮F�������u|�ã��������q4��Ȉ� O�nlob0DW-�h�����g�?n���3w=��}�^���|�ه?��S�~��}��~���0h�� ���Cc�9�t��=<���Fo{Ǔ�m��3�����holƲَ)��8QWb��)���{x�8>8�����1Xqs��?ĺL94P(Uoe�K�x��F��~�)��3Ni^�)��"n4D^,Fރ��E��o���*vi���{#XG��]G
���O|ng��^
�}�D��Sw~��O��J����p��6
�s����@�8`_;o ��g��&0���9�U�[\|~������ˀ��t�F�W�(�ρ`
����S���}��E�ԫ�m~ ��&d~�5�M�t~Q�$ӵ`�g��\�c.��FQp�h0�M���^q�x^D�����X ?>���)(��y���a�ts1��{-6��8���[�htZ��:�q�������������G�������������g�����]���w�x���o^}����q¼��ֱzp�a���!�~�h��1Y��g�v+ڣql�;�b�l�!��N?����r+�o>�YDZE����"�H�+6k4�NI$�)�!�)39� �����H�9 ��Dm�&���6*QB5bqx����'x�+��ޭ�|�6H�+�T�@�E���2��R��h�D��ύ#h��?Ú�e�W����n�T��<�'��`�8����%���[Id{g��k���k�H�u�)F)�����H��{���q~oT�������Ueb^��������\�K.��u�|����U	T�}L�+X�� H�n����c'J��eA-G �F�������P�L��o��M�͓��0"&Ѭ1Aq��*F�V�lm�hk㭡(�h�bY���\������p�G����x����9b�7@^����3�x�O|����3�~���k���^��m��j:���Nf��cY��<��\�k��z��F��ى�`\X����h�PP��	,��ڧ��#B݀E�肋nN�E>�R��2���k�Z�W:r�1��F�<g;��u��+�_';?)6���Y�����Kсc�{T��
��8���K�?���6\�?k���*HpL�����%0m���֮���_sM��w��I�(H��tK(���F��,���ug��ρ���=�N��  �k��a)�9s�l0����֏q����:�����#��בr�lܢ@�kfD��E]PiXT��x�[ʇ���t�‎$����8�ݏ��;���tu���a��:�f�ƁYt�����1���щ�3��7����bI�W?:���o�\������;���>�b�/���/�������>�K�}��_sr�fwz�+pl��L�b>��b2�$4�w�=2�iu�XAj�:�`1llFk;Z�Ml:Í��;��Y� �qX����V�/ �^U����97GWNAe�Q A)r�
�s��*3���l��7�<��۴W � ���1p�����	ʰ+ �#W�Ju݋6#������f�A��-���q[����FQ�2�9����`�{p,�t]*�xi,i(���^�/`P6��y�8�C.l�:W���Soi���&u|x�͇��mx6��4�����U��|n�O���>�5/��7`Le��G�ErL Y�G��I��.��z8�T��Z��d�:8��uR$�Tj�^���Ã�8څs܏��q4V����$:_��l�g�"��!��Ƹ㭍�6���D�3�vCs웽�;�����v������_��×@^��Gz�>��v������G��d��<�ϔz>�:����[ $ x'��L8ȵ�1c&��0e��������lmE�L���u�M����
�P�}�;�3g���frW-P/�P��p��Jt�b��Ǽ�:2*)���@-�rh�����������d>Ҝ�����Um^���Q�Sq�Y�~c/R����nځcv��4�����IYxA:=��|.�u�ڣ�ӂ��q�8�j�[ Ň��h��y��~��FV�,rL�,����s�|�4�Z�M��J�9D��N4ͩM���$I�k���i��ί"�g��{08
F.M$�<�׊�M��| �1�^�gTV�L^^<�rӣCq�'ǁQ�j2�f���+��$� 2��^C27�fWr豈v��zȍm00ﬂ�z��F'��n{��c��{�����=V�_��|I�O����'>��4ٽ��������I�&�1�˙�0��pµ��d^ׅ]���HC�q$?K�ѐ���@�5�����mnǜ(kو6���z։�U��>��H�V�9�mUb���S�,�$7��Ȉ�t���j�Y�iN�ģ7�]�pA��a�qYw^5���LBt�+_�NX<g1����$)],�BD5E㳚_��]�`Jϳ��U^4C�4�|Yj@�9|>�y���N���BR� ��U)�A���|�p|^c�@���.A�H�c�M���(Uf�xy~��H��E��q�YL���r1n. ��ye�|:�E�<�;��2���cpD���8�a?H�#�� :���&��h:��;�c~r3(.���h�kk�d<C���V��4��Yh��[]捷��1���3�5�>(���1�w�n��?]��5�k��m{/2�7y� �>���O?����ӏ����`<�s5�ǻQ�db6���V�&��/Wي%�&��8�Q(I�<�29 �Ԁ풫ъU�s"�� F�����Xvz1���?�_$�=��M��}������2�M��,����� �8�?:>Y�0�^�&G�|w�e��^���sΟ?�����X��?��Rn�K���wԼ0��6 ����bq\��cp��g"H"[�|�8��A�|W)��Ȓs��y���2�0�Kt#��í�Q�8�RD�9g�$)r�f��G����>>�)��6A�A�3Uk@R��G T
\N�Mg(�-�	�L�����P���q�[̣�R�/����bʂ�ǺH�#5�|�����3�z��R|�Z���(f���f� ˫-��R��J�w�6�e4�Y4���~�E���V�A^��6�3hk�"cPp�BD~0������·.|ɫ��[����Q�?�[���>s���ߺ���j?jǷc�3��z�.������v[�X��1�9�g    IDAT]�����M��	N:�1��]j,(Q$]4�f#��i��ފ�p������� c =`^`U�4/f�HE �4����q�����:;���N58~�_���� !�>{����}���@�*��X�4J�]�G��i��7�%* 3��DQ�A<_���;��T�ρ_d �Xy2f��R�R��f�hpT�W"J;����y ���J�"�"�����;d�..S����W�q�ʊ|�Ie<-?���I?c��9�<V�Q��Ku�D���G�cݖ��jZdB d���uoԳ�_E����{%7�T��繴�hr�@�yዙ�^��d]�A�����!��h s⺠f���A3x"�9��YtZ�yz��ׂ��:l�t�գ�^E�K�Њ��F��l�dq8�h�\9߫��|�?�M�顔\� _/�����������y���r����|?Z��l�cα�� r�d�vb�d<P=��;S��@�����uc�4B���R`;���!��ъ�h��F�_������16L6�qD�S��������ŃC�[��2gg錹=��R)/�T�����W���l��.�vJg�U�@��^�%|����k_��}�<��2����9��ӱ��Ve���q�8���D�|�uU�� �>��2���x��\�`�1G�b�St�st��Y��X���xc#���s���eiF[ w;���LO�y~Fji;g�ב-F��bp��H��h�<�k׮�Vϣ5��6U�t�`^V�!�)�5ڌ�Nӣ��Ȫ<7"]�b]���[Y�@r��ݤRO[��s�}�5���
+��IL���$M�q��=T�!���f���z��-f�<��t�~��1jnԗE6��E�����Z��n��3ތYzl�ht��y|�����p��K ��������}�3t���Y��=�?T�g�֎ƪ�E#fs�F6c!?�ڟt��J$���k�QðYW��
D<�A���}/�U��nG��z��~O ��WD"����0���/��d��+���VRT�)h�?\��fm���e���TIdxC+�"%T䅦/��	D�oli�3�������{Li6Bo��/�����*�e��W�S�g=�وÓc-*s����U�=Pd{^�[)c=UJۊ��òx/<���s�u��HN��^[���F�P�qDܼfJc:;+�l
���c��t�X�ҋnP�h��:'S�b��/�E�f����$�P#.�U9g���,��/f��䶳���fޛ�K�M�)��g�|-���g�|���}#p�kAM��S���:e�|<><Q��G��P%�T��*���W�ݢݑP���/��`�DԘ.��9����z���7Es���x�y���ݹ�����7���<�zz�����>O|�_��S������w���,��]x���2�+ �����EK�5���y�D��%����F+�g.�q��X�~aN o	��Ƥݍ��3i���Ĝ��A�$�%``>��$e%��U�P������z��C���b>�G��S���T��)�^sI��3�m�V�^+湜���7��ZHO=�T|�s����4��c�Iݼ�S�*��(֢�j�{x|������kW���
�ϟ�8==����@��	���K��)�|9H�Zc��ק��c�9SE�-wf@�ǽ�����3���ˉ\yM�ψfF�"H�� &�L�$�5�H�}��V���뗪��qV��#�J�x��s�	�M]�|�*�Y���=��\^۶g����R��x/�~bzp��.r:	L�������x* l7�1�i,E�A�Y�(3E�<yN��@�l4W� %gY�]�IF�h���]��G�zٟ�o}�3/n�$ �_�W��G�o�<��[��Dcq ���8>blE}��V] ��g� ��W]�n1v�D��*��dF(]�?HPNg��t�����(�nh2:�";�s����0+M�L��y꺢�O� ���q����U��n����Sne�.�|Y\\�I��!����Ԉ�|IO+�e�/���ޫ㦒�(�,J���V]@p4Y����#�_-U�R4X)r8��^3u��Ma�-�际����f]K /Ƽ�S/n��)$����k�v�3��)��^9��"ͩA`�����!��^�`�X̦ٽT���5v�+���]�g;��AaG�b'+�v
�&e�t�@�xG��0���B�^�+�x��\N���X�Z{#vu����Z͈ W2�8a����6׺|��Q��zT�9�?;���ΧJ��2YNu)j4p���Q�o����*jp��Z4�A>ފ�x'v�y�O�y٫����G.}Q�/��?{�����j���k_��t?j��Tވڢ+
3K������%@�dAJA���0��CZ��+����W5��hw緶��}&ڃ�"��j�'s�_G�VԮ]f�8:ZKrX�~+�s���Im�5�*y��0��Ul���;D��$��A��L��^OL~����ʻSW�9s�k1�d�N{�qc���b����DEN#O�s�6G-�Ʃ���ڑ��㪀g�Ͻ�N-��-��E�%���ϔ��������h��< D~�^X��_q����qU��uf=��E�mO�zQ!T_�Z�!�}��7!��ˈ:i
o@kiN9>��ܴ�����s������}^2��L��\W��$�X׋@}>9�;]1s6�C$w��)5[	c��1�;3��+�D���av����o�z�~��4j�e�u$��,5������u6v��}��w���?�~���@�¿|�����ݿ�:������h��dc%��U;S�9�uC �$�T�MT�~�D�k^k���1���f��fZ�MM�9ȃ�	f
3s��S;"z���V;'� �^/��b`b`�?7JU��D���k�}'A�ǸW�c�E~��YKYT�V�J.dG��K��i�8(:4�6�.Y�����뒟�©T�����`���8`���$.�'?K�M_sIEUHp���D�4{�ss�<[N4`�w�ꨨ6�)R)��T�1��v~v1L�1(��=��H�q�)&�X�?��s��H�E����kZޔꄜ���4�:�
���~�y|0�5\�rPJ>���zP܌DoT,�pN���*��4續x�=8�i�z|����N�oĦ������I�����X��#�� e L�(����s Ūk*��xQ �\Q#��I�汬%@���h���aWx&ν������^�_}��������?�w�3����ɳ�	���%eьP� IzMt�E������r׈U��IAJ9�!��&���0�'�9D2)y[��v/��P��-���8���c�EJ�L��VG�(�P���D���'��rB�'67�v���bqT����@�d�REVƤ��w��"�i՛1_1����a��CmW�\Q�c�zCr>��{+�*�g�R����4��tf�w.���苟�8@z�k3l��������:�Yc>[u	�Y-���Q���m��o�����S+�.�� 2��������H� |1�p�BU�uf$��Wݸ�f�é)�H�e<L�"�1%��$M,�K�����\�h��ë�Ո&���D�\���u�1[*��d5z�|�G�^��0�S�h�U�9Ʉ� �|)����lu4��Rh�x�aD�M�q�?E�� HJ��G�B(D�lx1��X��F��R=Ꝇ�Z��8��W���|ݻ���?��U�S���}�_�������6��	 %:�b�`����R$9[42}�â���͓BLG�G|�� ˮK��Z���_�Փ��Pm��X6Z��_��uK�Y/"�f�t\�s�P{&H�4�Jm���ujX�8E7'V]<�. UV�?�#�t~����C��\�h��#E���/���P+�#Z ��$�.i�9U1�Q�7z|t�L�+ �E�#+��x�ɉK	����� ^k
@��Ŭ�(�/�KX��������U�c$R)ql.^B���l���M:����^"�C�תKv�UQV���y.L�V�Og9��g�> <Iu�a�L�Dw�
r:ěvpJ������L)d3Fب� ���������t�,DE�~���Q��yQ[?�,|��1q�XȈ�矧d��#���a<H�K%���huB�2��X����G��C���Z�J��Bo�Cr�门 � ȶ"ȝ8��~���_������|��
 ?��}�/��?���ɵ�ע�<�e����A�M�Hez�Lӂ�H
�GV�>��
�ي�l�Y�,`�,��)��;q��ȈX�T����5�1#"�Zf(�uSf��B"ήg!F2��v�9Ӱ2_��q��*b��4�첅T���s1՜�S�ɩ#6��C��rn7d|��T;AY���MNū yM��q~0:-�`�긋E��>�j��>��6b^��P����P$AE��I�&���"��k�9���eu��Q�>ޑ��a���q A��B�^�-w<���E��,�*�_�鼸[5������x�]��y��)6R��ӹF��g=�v҈��Eߜ9�X �ʉ��
H�U\��s�W\�W�L�g�U�f�<�`�{6���%u^���������D�3� �U(�� ��@�`-�eF�r�2f��C�}1���\�x>�4<��M�M���s�$Ҡ�@Z���N�����������+_T �/�����~��~pw^љ܊��Q��j���R�&�%�#B��\��"b��H�[��Xk� �G�pJ���1�Q���xJ�����R�X�a�.'ppL �7�J� �4�2s��m���T�Y �x=J~L�Q4p	(�.�ک~P�/�Ӏ{n"�vd1�@I��q�~��)91"��t�<��2�~�Aޜќ��c����_���MY���R�_���<�Me���S�����)��Z$zX��ہa�`0*)yN"�:�?JX���8�LGU��"��g̍0���b=d+?g��j����:�UV����I�Iq�{�stj)��%��<����I��h�bS�K�%R�f��\,<=|!79�#_J�K�%��bF��Lb�Wr��/�P-��&�Sd�͂XQ��Ԑ1�ܻ��Z�g�R�o:��*Ҙ��l��{��߹��|��������/�����r����؜D�V�ԴS5�D�� �ֱ��.�������P���}K��l�7̒V,���#��!%�����7gw��A=�N���>{$2Ȓ7˛SQ �C�X���G
T�OG�ML��hs�e5��:5��~���yi�^�:�����1�Vzn)���Jd?��,�X��"��k��Aٸ���%90�Z���N�$j	�u�,�qq>�2=�ב����,�^�ˉ���ܹ�[C�j����s�݆�x�]&ހ�)hrc������{��R�2G��K�La�Bn*��@�;�>��R�D8���=�������,@�u�ߖ%���6`O��К/�ȼ�C����;�b ��t8#�,�8�V����ɀ>��I���z��KY���\ YG�yE��GcDG�v�������^���;���}q� ������|����ۯ  듽\vS�dve p)�bsFE����38F\|H��/���\TI|$�S��"A�h��F͛T�]W��U�m?V^�%��s�۲Dx)ա���<e�����Ĕ-����޴���ҋ�4�ˈ�J���'?j �w�k���!/�";> 	`��G����v>���x9���z�Ze��!&����t�N#
Ig�"
@J@�7��Z�� ���X���t5[=�!4;:�5���R�ը^�6_ތT|+_>��Դ�����"�R7��Q=��
�9.�t�  ���_�
���k��Ɣ�WRLm�AP#�A9<�Wf�4I�Op�u��Z��K���K�+%B��0;w���L��-�"H$ŗ����H�>m"IT
��C��[h��bw{Q�=:w?��e�|ݟ��ȟ��?��|���:�����"������_��3H����i^��̪,_�զ�M�x�FH�v��e0VڥVZiJ?�
�6biD�toC� .	��#a8 �鞙���K�Sqν����j��DD�1�U���;߽�{n��B�����[�f'$���_-�$h�΂Kd�%9.*� �YP� �*�	�,ژ<CS7&�Q�z�����#�ɇ0Y:��!T{��F�����2s�!��>�O�q<
W��?2"�ќ줰�O�x `Q�F�ۀ0����y5�L���)9G�ZL����ѐ�*Yd1����M^�$F�����4�U�r`�J��-~�c#[D�M�&�̌x��$�BF��詅4r��v����G� ` _���LgԂ8�t����]�o�T���6�|�b�严�o;��8r5!$_��O��G&9�F��;f�'�ױ�Dg"�g��񂢎,ו	�AͰs����S"
�M�t����I4E恹�]���7[99!7�&*�t�̇N��٧��7��H�����N�/|����է���Ak�T��G���A�s���&��1� D�	VC��o�!@�R ���4#��F�޼��+�� �֡.P��X����>�W��ӗ(W�5����uB�f�y���zls��I�HNT�½I�P%�4׃�l�wtb���l���{Ap�b$e����L�!"mp�y�u �F���Xv ��&8]��@AD�A�!�Ӎs���a4��Q�,�� ���% ���K��1�'D+�	{�p9�?�HHQ�z���^���;[G��ڹK�RZ�u�vQ��i��q��7W�+2L\�(ԋ)�*�LGf� ���T�D�,���:�oMSj���\�r�\o �H�� p���n�Sl?(@�S�ǨC���r d
����W����,�����3��O>�S�h���' �����鏾?�X?��K�]#@���I@@�� ŗ!"H�Q@녭���~iؠ�p��M�3��������"Mt�pt������E�`��{H.N�N�\M�T7�W��E� h��; ں8�wpo^�@j
`C��mUc3�A�RH7�{��E	
>��t#(ҏA�pPn&kt���S�����&��D�����o0�>��V�����,�@C��)� J��v/����,*���C�H�F8P&c���X�7O�r�yɟ7�F�s� hzO �v+i'��B�Ş��I��:i��#��u�7����Uk��aQ��#�\��Ƹ�]��R) 3�ü��?]%R����'���IJ�\�H���k� ���$�u3S&�9�T
�u��u�Uk�W� !�( $t�%�N��O���G�<��O��'v��Qc���' �s{������� �b�&�nC��J �H A�d��!::�j"�����:4�ij��E#�;R���:����cl�$���kDs*��3*G��>��L0��X[��a�Ũh.�X2HDnO�ϭ4��/ntf��W���[��)�v8��6����կR9:ߨ� �c�Y=V�Ҳ	�����DQ�!��������ϥ�!R 3`�� ���b�p��I7�VH��������Ն$,�{���<^�}�gp�@�5�>e+q�4��lA�o�J�ԟ4<,��:��:S['�> I)�ᇞt�eV��)#b ��J�2`u���B^���Ae<"߯�a�����E�!H�cxru�Z%��v{׏�C�A���1��>��V"�����:�RYr�����{e��C�yW����?�����7%�oʈ6�q�v槵 �
K�9���D�=��H|0��Qe.p:ѓP%N�{��eә�($��H2��q�����g$�p���b'*�I�\���u�kԉ�G/��~�$��$�`r��Q�4��,���ؐ�N�rQ�Z{N���A����R~��E�윍��5z�>F~f����.���0���G�L�b�=-�����dQ�I���8e�r&s�Ea��h    IDAT �AR��8P���:=�Y<C�k��v�:���^�*�`�%^�j��ĬZ��T���_����#MO~B֤�'�	��Y֔�-���I��^���ũme����D�>:�������"h���D�@���ܻg��jܱȼH�H�c1X�h@b�H�BC�0�? H��c���2;57X:~��>���x���]�>����� .@ѿ������Ʃ��&�V��o�S��F*�V1r�� !�uVЄ�<$E݂��V������.�(祒��hc�i;m�s�i �i�ú	��~?ǿ���b�#m�$ !���	�#�ѹ��V{��b�C�)���4���(��")�ru����)� �n�6�:@���0j�ע�f�]z��<��}�4 ��F��b~�[)ig)��� Κa+$���D�����Bjt���Z��G�\��1� �EG�`��-�$����{�d����U�������wX-���K3z?t�L�����שR�4�C@�y<h+�W.�I(X���Ѵ�ڏ��X�E4��8�w����^��g�8,��B�%�^bt$�˄�R�tڇ���4��KcD�I��0��H�2)����r��o���W�:���?|Ǔ��?~��q�8lȨS�sg�My�$�0�p��=Br�ߣ��+�Z}FJ�^{�Z�9���B�b������~	i$7��я"h�v�H�M#F[�\,VP�'ˌ\�B���n� C��B���9?#i����`|�p�D���ʎ*�01�E��)��K���^�����$#/�^�6�1�k��<�fr��r��lHx��H��4z$���¿3����x� �7�fd�m��!��l5�#&\Rw?Ҫ혟GX����3�JGL'\��)�s�8�`3w�d����e@��1:�#Z�r��~�D}����f>�(�o[:|�א6�"i�&?dL��k��+D�,�P{����D9Q ��,��2$xE*W�������2L�%[�����rx���O���w@~����/}�c�o��@�zJ|�/�R�.6P#��B	%=<���E~Ѥ=�d8a��(Ҭ��ӛ���fD{><	}��BS�<��x:-�(�����VHwd|�1�&�f�$ދ��|�t�i��.ε�S/V�L�M�j��v�(G��O57���W<-*���`h�A>ɸF\{S&k���]�:Y�F룶�������GY�}ԁ�!��ƊD���=��U��1��ݧ��mC�<���m�$�-�Ĺ3��GR���k�{aZJ��
V��5s-��v�J������?f�Ʃ�l"Jw���@2�G��'X��g6*��m�G�~o�}y�ž!dt������i�j3�6n؋:c�D[���ة)����њ���I�V*21�4�9|�w��>��w�W������`��u2ӯJ�SW�GEܘ��!o��Rc5����z�߱�ԭ�e��4sM\�&A����ɳ����k����&	�tu�)�O�39��"�FT�b�'�������"��
�����Ҡ�FyZj�E�T�l���BL�T�Ǎb���!j�tׁ$�뼝�$(z=�*����<������9x0�4�4�k#��|:�^�I��� t�_ ���^��{��-
��}r�M���r���q��F�a�g�k����[bm����b(pn�gCU��
 3���������C��g~��MD(N��[č��`<#�A����w:�X~v��^`�A�U���x��ф��0$��{�E�����K<�"�M�2��2&äH��{)�/�VN����{�u����������D����?��˟������d{W���aJ�C�O�;bC`C��bl����
��9TPr����i�N�qV�t��� _Z�h��zI{-ڠP�2�4��#�b`��[�QvgR�1���?O��n��ܘ��5�f�h�_��i���V���[�{����sE�H�+�Q0�:"'��ݒ�h�p��	�c�WnL�m�I��+î��o?T��x(cq�B�~V.-F����I�C��ֺ��ڳ��Ub��;.���5����)�< h>��Q�1�l:�kG�L-�y� �@
��~����K��{4�����1��{��n�{º�3��G$?~x0"G ��%�ǁ���:�5B�Sm��{B����,Mw%Cdh�ŨX��2�d�0k;�ץ�d'��0;?�]9���g���� ?���z������;ǂ֎$zmC�(�=��^X���n>aZg-��d��.�0j�+�����1�|F� A�*��!���K��I
��x���|5�Gc�qaћ	ѹy\�1�ӜȆ�M�c?�T�F~�VO�Ie�;���3����D�}�&���0��s�0�rt
�Q��oʟ��;r���>Sm�x���a�FRW%<�z��8�jkk��Fy�5/�D��(��s3]= �m^kرA\k��_^IH��Q�OAM)�p��OP�"m��c3����0�RgO����T ������N!�t��
<����)�H��`�:�;3�Wz0��v����C�,�
��Y���D��4Eڨ����X=5g�n@�+
��t�Z3q���� ���ʒ�^�=�G��������/���>��'ޝ��I�w%t	����Hy���d����lt�P����׬lG �'.���=�7��7�̉"�x�;�M.�>�𤡅� R�H����N5��#s���c�cz>ҧ�^c���a���v�dTH�^MM¯Ȍ<�)�Y�y﬒��y��)����B��7�/��%tM�l��\y'�Tw��0�#H��y�KX�}Į^P.Q �-��:5����f>λ���k?��:�\��:8`8H�@1��#i���gr`p*���H�o�������X��n
ߋ��D}��F� ��<Iu�c��@N�v��5o�S�>��"�'x�SG�z���U�i���i=+�@����$�h<<�����$f�8@j��	1���qɕ'�(���g�������]���_��g>��wg{�+A{W�C���ׂ[4ҙ8RME4B�VB��ָ�QZ��m�y�M,�x�rlH���	J���n�����c �Ԝ�*�>� �<"waD�4���:���0G][HPBt0�~-�}����.M��w��7�[c)Oq�P��q�BG7���l���d�Yb���98�� X�穄0�L��;�;��3x����P�d�Xlb5�0n�7�8��Q#��(��O�=*���v{�E�(@�P�<զ��2+� d�kck=��u�'�X a^��i���
9����4�NEx��,����[R�J�$�4�wV����#Jw��H��_�*�<�kt#�H�:�����Ҫs��I���Щ��@�&ތ3htǪ���z�a�|iBⅢ�ʳÙ#'�q�������6����7 ��I46e�u�JJ��4��W�.��Tǝ{�p��	�"� ���ݡj�(fA�{��^h� �K�R�{E:H�H����KT(RW�Wa����G�Y����n"͏x���	�M|G�/d]9���*�G�2:K�ٱ�{��C�u�cA��ra:� e�5����G-����7�'��q��;f�
��ƫµ��m0��~܉���ۆ�po�a/=6�kG����p@bU5�1��a:?��Y8@r3`��m��6������:L�=�(�魲�&*��8G��X����f;,�x7���94R��!�����L���
3�pՁU�/ڟ�iX�pHF�WF�֊�T���wP�H�tJf� 3@����7�#6b���Nјb�
;8|4ch��N���G2
�ḅ��fGӇ������?���e�����z�ן��{���C�^C�a�=��X
�0t�!z��b�+:Y!j�V�$�Z�m�g��Lo�K�M_:t�qZ��A�Z�r���_�Z5RDK�F}���i
�H-����ø)nT��H�"`O�ؙa�����Bݢe�9�1� ����=�{�.un���+����۹9�pÇ�������t�D�j��1)u�9L�\Am�9f��%1	2ʽ� ��3�߫N��r�`
�=틈��s� M�5���1��O�R��nH���+�n�I��A�,a<��ɨ>�}7�e�r|�E#[@�p�2ݢ=_ȡF�L~~�{#@Ĩ¯��1~������O�΄���i4��z�:@�o��."C 9
7�����j��_��1�Y6���KeINLHnrF�+��q��]���������'��o,g{UI��4�@%{Їf,)q�}ԩ �vBVO�m ���zk�4I���r���F ���j�5�%b![��cO��ճ��6�1@(��Y�Hwzr)������=
�(<��t!܀�U�H[ �H�̴�0�Cl������ţmFQm%�]\K; t���L�i! ����n�(Yw��H�Z�=�F\���@V�a�̢}i !"V����RmDѯ��*�_��w��$��)��r�t�3�������N��+�"�񀳋T(���m���N?��#q�{
�{ȃ)�FI�@����0Ȩ��]s�qԺ�<w�<p�
�V��% "Cl��cn��Y �!�/5̂i�@2 с�QCon?!R(�AfK3R^:���3�����_o�v��������|�����g>���$��Aw_�^�:Hj�0�S����ׅy.��a4("s Wj���U$���VSo�0��
�)�s�Gy@Z[G�U��A���F��'�<�f�������L#��(��^�H��x^��kq����������9���w��^�q5}���UTO;�h���R߼A�b��;_�+��숀:��yX#]��{<�~h��6!��g1޺�nFPѪ�r�v� ait��p�� ��C��j-׋���� �ך��H�Q��$i���\qW�� ����v��_��:��ꟍ6dgs�&m�#t�@HrށeC�x=X\Q(��4|~�@�b�	� ��8����3@��� �L� ��)�OΌ*ˇ߹t���/�~�#�z۳���77���=	zH��v��"��U!��nˆvxh�O�^�Y}F�T�,;2�ڨ��29� ��U�pC)ف�7���ss��5=ڡ��	�JFN_>���%��`��GHa4� ��HE5���!J}9`(7��4~��qP>W���H��Q�n�0��pq|V{.O�y����f���1�a�""t`czq�a4d)�?�kL�3E��yu����|޵F��X� q ��]�wl�s�;^�2�m���G���w�9��# ���Q.�F��2����ϩ�i��N�-rt�:ތ�z]W~��ß�1��E��,��K�>�M�t&�M�\�� |M0ò�:�ip�
Z����g�P,�&�b4zE��K�,���s��$��1�i�w�qIcht�S����w,{��:�鏼�G���O�'��\Jw�$�kr#�3��-�[ݯQ5��S2�����z(���C��=��@=��<���e�� -���hb1��4���،A���Nݣ�F�|�sw��d��`�4;����<e�#`|>Q���
�C�ba�� ����Х!	�@]�[�!��O� �X�z�� O�y  zIC`,� �`��("��# ZF�x=�ֳ@��R�o M��r�WD���Y�*|�n��f��Z-Z�^ϰhR"��SS/jX��Ag�+k����U: ���S�1�Y��$;�L��@HH���SA���������A�B-��;+�6�3�M����'ӿ��'�«Ξ��g���0���D�ǔ�� �"M�\�lyz8�x�]�G����~�_n�1�����H����������77��I�;\�:�;5I��H 	~ctr!Sjh� $� �JYe3H�7�piC�j��A��Q>O��{�"7Ǉbv��d�l
��Z���psX��vOًk�-ѡF���7�Ȥ;?�ى���n�r�9�2����\��m��==0��ިsd^��u�vK#!TR�Nm�	���
����S:�4�����R�7pr�!;�0:@��8<\j�,�F�Ӽ��#.��� Cp���IEP��sn�A�[�T�:��^����Y�>�ѦMr�"ٝ ��I�B�nF�A+"5���B���k�2/z<���vPh��k�?�e��J���ژ�P��.ҕ���6�D�!��[N[dG��S��ry������ۧϜ��7�mvg���~���ޗjn/�;9h	��G�� ��F2��\d����L75���z�{7�C��"�Cd���a��;�;O�X�A����*6O`�eX�xO}3��bF�(Q'�� �iN`�-����h��E�'�ql�G�L@ ǃ����g�@�`b4a�M�&i_#23���)��i��|�;�n(3agt��j���zSM�\���� j�A;7H��-�%?^	�V�� ]&6=�����kbl
���P����x3���1��X	Q�a���Q'�RI��~x���IYT�ѐ��6;�t̬H��*HJV{P=DF>x�=�d.��.Gf �y��7�,��Ǌ�Pe��\/G�Ȉ��7?�\��q�e�<��q����*��"چt�-�a����"bԠ@#IS��K�5}<-�Ce<p&M�\�̧?s���,��������~�;Z����B���y���m_���ޟlo.�U�u�����a4��*5MsQ�@��pD�0����[��і�B�̍+��G#F@X|�E���|��2i_p�_���P���E<6�^����d{{W��A��3�:Z�0k�F���gsC��D@j��jբ���ͣb	p$��2��"�A[��Ya�IDOC��	�8�{v�h$�0��D鴺ɰJo�7akB��q囓#<|�I�F��,2�	�d��KjC��) ��^� ��%��@Sb2��Ld���H:$��Rބ� ()��TE�-1���:��\L�ڭ�y�{��ū@1�{7U���GkH9�`����X`�ŸC�����_8���&��ӵ.۪H���HdP\�J��t}��0t�%Pu��N#0ۈ�wS-@���	����A@ m#"��PR0���C�����X��u��{Z��������~�S�@��I�=橸$�	Je��^L-����_��O=�����p�{"�~������~���O47�`�������1r��PFЎcP�b��&�!(r��b	#Pǈ�Y��.���
��o!�~-�k2!(
�x�Dn,pBMH�ۓ6wN>�ݛ���ӆQm�tf�F�*�G
��:���ztqn��px�"�����wy��w���w�J�"�z�R�p#��>#n< Ցmp5$�5��<�+Z�H�"2ي�3F���  �lk��Rl���c&)�l>t0z��BAJ7�4��?��xx�9��ÆD�륇)�.��I�#���c����^i���i��"�4�5Y%GČ�Ɗ7ތ�B�K�8ͅH��]��~uW1���AI��!J��Y�9J
7�WE3�$@]Mky���wW�P�`�W#T���C{��#��K�f[#k!�Yi�Q�-�ι���&�H��7:@R����n8�LSo��H��a�H'$��Kr�$�����ұ�:}�_z�[�27��~�o��_|�R�u �4	�4G��cz��n`�xWK�p��fp�� � -e@tQ������2�l!�Ņ��"F$�b��f$���l�91]�hx?�.0�u�ҥ�d �vGrق�Zh�ה#a�9,.��X4��rll,���|���h�)�܁"wңV��4�Um�6���G.|�0c�T8@�\F����`Z�<�Q�-I�Yw�a���4,�CKU�k�ǁP�g ��Dd��Ub����4_���?�2a���a}��[C^圱�ɹ���vgFpS+    IDAT������4����Z
��J ��p�Ļu\��I�ؔC����Q ށb}����N5P7J����t�;"O�]F�pI��H!?˸�F�IT�M
�/"D�=�_E�	F��n�hd���"��u\�F��V�{LCB7�K���
�f`����Q?��� �hc9����d3jF:�+�� ��䨴x�?�<��/�u�>�{o��?�{���+����F-�5  ���l�L��N ��^BzH���� 7HF�0�P
M��?�67Sx����H4���3���&���A6�98�|A�񄴑���h����H���ۍ����V9� ���eR�0�胋�[z[�>��;ܯQ��K�D�}��~�&SA��}@�p8����~�I]�3t֘��x\�G��>w����X���1 D���e����T\R��r9ƺ0'�|
��3���� @!8 �C��f�xax?�Is|�IbF�=�CF����{��gno���~�����Ko�7��S��t�1š �]Ua�m�o>��!����2�5�JY�Ɓ��J"�1�>av1�K&��M�Gt�TȐT���I��ZI�|ʧr\�.$�d����(E�5`��0�D�@�'hEŚ�c�l �ځ�C>�Q��k��5f��
�ciJ��&� ���TJ�e)�.����w~������֋M���?������l�@�!"H]�l�Y."7��a��Is���fg4z��N@� ��j�7�ܨ�!!}I�!�II�P�t� �Ҕ��yr �����I�c�#�ܯV�����9)�4G1��ؒV����i�8t	�TT�i1S7�X㔍��;i���p~�{ڧ��j9숺2��!.�-�ѹ���Q;�y,�ei�� ��H\��9W�t�=��0 �P����D���( �j��L��֨�%$@H��iQ��$"�@��47m���a�^�^G92m�TW�`_iz���� �j0�7H�<W��΋0��� ^*�d���A����[b��ſ�@�]�I�����'C���m�hV|����'#�s^�G�~k3D*�e!|z:��t.+�L��9�MfUv�=��.�s�ђZ�)�zK���:�:m�� �uH��=�w��%{ZX�)
:I�zE��5%r���i0d�=Ŏ���{��ݙL.}ߩ�w]'�g?�����_�ɇb����@��8]T�BL_h��� bc���
���*����$�Ά�;�������S1���R���d�"�ʜ��2�Df��66#*�̡B��QhL��4�-:�T�SR�5�)�ڵr��%�ԥ�nK�&�f[zݎ��Hױ��Y
vЄ#̲���(8:@<5>VR�8�)����jأ=�k44ë7���Z#=T^q ��t��p�NH��b �7�'$]$�F�ݓޠKNY��#L�$��JR9Ie�d�Pϋ����5?�A���I��~��`ĸ�w@Ji")T�)&��8d'vm�Ѓރn����W�],�G�p�Z�E�; �@��6a���ot�O��?��4��0�e4��r��I��5/6�L.M`�����:zQ&��uE�+%��)�� �"u��f�7O�0r��7�Z�!PB�@����� �vK�ͦ��m�e��|	fz�7�V����kaF]Z}���
PJA���ŵ�$����grN�+�������o�Wk�S�����"�_��?������%�[��aU⽆@歄1W���!NF�|�j0��t�vj2Ŷ�i ���g�}iTى���������dOd���p�tr�Sx�����r---���<�r�,���r��-��� k��Y`���6[ҨV��hjU���h��"�G(4�ts�qD�i��Q�$w	���7�W��π!��_��w�N���3B�3��m��C�֋�8`,@�����.�	��$��rl�xH&?)�lAbɜ��9I���HP�Nx^�?�ݢ������,���e�9�r�\�tIv6���S8m� a/��I�׍���ڔE�vX�J���bH
z��]�K��2������݈֨��<����h��c.��~W#�@M�t5�O�D��Kr�q8�%_,J�P&��Y Kgr�Q�ᓵ#p�!A#�Ð�Y�`��R,N���lln��+Wdgk��t�Ԫ��<�I�ļ� J��Ԇ�
�X�LH�ՍRҠ�M	7qH��2�x� �ҴL,���釞�?�:�|����Ͼ��?yO��=��vMO�D@pt��m̩�HWTC�҅0���r��uX�H��K
sg� �J4��I�LOKe~Z�-J�R�X�V�()����҆0�zL7�j5dsc���2U���쬬:B���ؐO~�r��MF2�z����j���T�w���������bz:�Ϲ�S�+�ΙQ�A3��*b�mam)[�
�E���sY ��o3��L#*�+	�JMP�ژ�%%�OK2�01�."pO���J�219#��9I�s���_.%�T���r�.�ͅL2!�
2�/��������ψ�dnnN��V��ի�կ~Uοt� K�4�R�F�5axm�PU�p�ޅ�`��e������P�n�U#�gQ� �h��� J״�[�,��I�A 0��{�z�t���Ҥ"��I�����Č$Ri���TZ���mi�����N��:i���	^?\땣XӇ��_z�%Y�y�3n�^�oo����o�Jn\wp��5��$)�?S3@��������ޑѳ�V���$). d~jN&}�䃏��]���(����'��?W�ڙIw�%5�EFڥ�G:�m4r�@�Y����5�u��b"9�gY���w�����dYf���grnFR�E�O���t�P�g%d��;��T�*w�L�k��lԤլ3�>�z\���>tH�[ej���駟���-��ޖf��E�D\jU���"7��Ac?�
ؤX\J�C�~R����m��a��\��R��#�d"mQ
R0<�OMt �4�}�����"���y��*L���H��OII!��D��^��E��P��|iRҩ��*�R*WD�JS4�Bd��M��k��FB ād�^��0:���f1�����Ԕ�=s���+���%^y�Q$$ʜ��!��t�'#P4ب�dA.am��>r�<H#X���rs���lp!���������E��2��S�**�&�i?��z�=�K:oφ$�	��S�7 ��b�$�NW
33��S�Y)��$���8nL,`��3�Z�!�6xr5�@�]($KK����].N��aOO���<$��\�yM^|�E�q�:�8�LJz�������#�;R�֨m���3�dh��B��j;�1�dʍ@Ҳ�5F��(�;�G���L,,��{�����?s�X����<�&@~�?�������4:i��`��P6�VCt�`����0�H/H�M��n-� �f"zΉ4{I�r��S�zꤔ&�2i�1�b�<�@��A�I��V�K�V�z�&ս}�vڒ�ܤ���ey��>|X*�s�H�?���L�������n���m7�n��p�AV�'Ջ���	�Q�f7�@��4� ����ٜ�@�6�4����vDhT�h��v_�j�E�ʙ!E�C�˧YE��;e�R�TVE���H~bR
���$��$S9ޯl�Hn,[��V��1�V��C����;��8$�$�Ͳ0���ȑc�0����3�����ҋ���΃�]��:�ۘ�7�A���B���>ui�`�~��H�\#�����TAoQ����8x�1"ķ���н�&4�0�%z�9�[Sq�#j&UR�!Z��`"�o>�l1-A���@�%W������t6'�\I�Ų��Y��F,�T�u��j\sx]d �l� ����e����$#vPY�3�\Ӈ��0-��kr��5�r��ԫ{,8������W���m�Z[���}�ے`��r���8�=���@��M%b}F�Y�J��2U(J�iqR
3��<��k���g���� �A��w��Ͽ��O�7�ݝa�!�!�A���s�LlV�y�������h&Mih�2�,��!z|�I���J�e��a9�������b�~�),�,*�	�#*\�K������r��{;4����%��T�R��������8�덆|��'�o^ӈ Q��>7�4�9�ޖZ�*�Z[z���G: L�)��ks��Y�͙V�F�X��r1r�4d�d�j�m}�qVt��$Ɩ�*��W�*y C�K&��T6.�rV�H��)M�J�� ����D"'�\Iꍖ�2 K-@r���=�Q�����>�*����l6ean��4��&&�2?�(G��Ƶ��o>+�Ν�!�M���Vݗv��M����^�U��ii�@�,&�� ��� �#H���p��Qc������y���F��;W� �sc,(K�r	p�(�t%�KHy�,���%���KizN������2��J
�������_�k�����Y���;Z��¢v�HB�=*Ǐ�� �R��e{kK.^|U���Y��l�v��z��M�q�4�2��FL��;(�cc_i�� O ��� �?��� �x./�|^R�����#����'��w@~�����o}��ߟ��Ϧ��t�r"��ƀ�kl�+vu�mј8F�
�MLH'�*􍩔�8> KG��ʽZo�A�%Mp�XF�����Fv�^o����j:Q(Ji��E535-��s����Pp�o���7���\�|��DZ�z�|�vSS�N�ΈggsG�U����Ht��<�Q��C��6��3_Gv��_ �xu���\��>3)66��`08�qi��)*}I�6����EѠP���Ԅ��}ɗ'd
vjNb��4; ޳R(NI&���8[(2R��R�plkfoEH%���*�#h���eI�2�H��9...I!_�aYo���oC����I6��un"���cʾ��#]\sD�v]IBXβ�2��dTm��{l��\O�'�
��1��:>l��F����Fvp!�S1��>�7Aw����8��ə2�Zh[��'�;��ȡ �x u�1ʦ�b��~Ԝ�!��a����5�WbM��K2�h2�C�}qnQVW��te^����l=Y�ܐ˗/���&�g4I�D��3��w��浫�&��{�:�(��
���D �h&�Unv�$Ԭ#�J�C�@7�d.'	T�楼��G������8H,�O����[�����m dU���@r��V
F�` �֙4  D�(�Ж���6N�K��Cr������3����f�-k[[�����A�%���cꑟ(r�4MF1���'b<��cGV�����d)�iv[r��U�x���z�.�z�@�Tۇ�mV� �і��=�%��A[�2H( ,�b�(���R{V����yo�s)60�Q#�VO�њ��.����g�*��c������Ӿ�Ԅ��MQ��gdvyQ&g��l&�FWm��e��/K������%�j Y�U����U d��&�냔��di��5"&�|��
�%.;��������]�(�%�N3���� "��ݖ��]�[��n�%�VW����2�cuٹ\���z��i\�`I+�А�vWq�� �6��D&�2����U*ȣ����Y�](Kq� A.%�Vdn����ɗ�������o��Cj� �En�Y���������T�"{�����������������&rk{�L:�{0�L<%�T �vO���x mߺ%۷֥�hH���<
9Br����)h�.;g����l��n�tyV��<q����?�/7���yǏ���z_��?����|�r�n�k�t�V4t�8@rhW")=�d��ĳY�k6�1��Ғ�}�Q���ǥ��(�\Vjݮ\�rU^�x�)4@�M��fԊaC�>`�2-6�D�>���}�> �B����M�!�/��d@miw�L��n�^U4#��w;L�H��3;8 H E�׸��ND�&�@��
+�C��`�=�ݟ�3C��c�Ulnl�05t�-�H99�HD5jM��R�,��\EJ�e9|bU*���@Z�ڗ�ZS��A�6uA2�b �/��>&�����5|���@�0��k�͊�q�W&���R��f�6����\��������ѱ�T/��
� (�[M���zUv�dw���X�Q�l2&O�-Rw�l�4��nM�F@�p\#o�$}�$|F5�4cf��C�sڡ)�H�������,V�<S"-�t���e��kJ�֓ť�R���������4S!���n֚����v��b{�k�(������aYY>D�D�N#iB�Ȕ��=�t�ܸvUڝ�dR���|�ZL�]�:�k�dsS֮\���5���ɨ�&9��{�#܆�Zؕ�2ԥ�0/T�9�'@�aFż�G����<��c?w�u�<��������S���dk_b��$�����ܔa�#��HA�X�)AG&-k{�T��{�<������`��i7��\�qSn޼)ͽ�U����쨛�e0��ەV�+A2%�B^r�#"Hz|�a�$n~l��^�͝MF`��bi!]���ը��y���dU�_�Μ�=r��V�@Y?�J�ޔ4�H~8�A�
L}�"S�Q��z��zk��cY��F��ʧ�02�|h�������" ���dQ*3eY9�$K�W���{d�H�n�&�[���$�~kk.;�rT&'+r��ei4�jz �����.;����$�!���'�W8�ʡC�ea�����
�AWtG��qK6�����5rm�*�}vz @S xؕ���Ei�#[�r��5r�8i;��@tOұ�AK����P�p���-��x���;H���#*õ�=@1�l��ɣi$�JIf�&	�K��ȩ��OH{����i4�2;�̃��h˅����X0����u���(xo��i����,��ؓ�=���գ��x|h<%uhTCj6�6dks]��]Σ	b1ɦ3���Hq�j����r��E��ܒA�����4%Nc�aD���� �,�N��*OHqvy0uh�O�~�/?��ع�"��~�=oy�KO8��]��wxAG�X�%�mՀ-\���Y�D�ͱp-��)uhGH��۵�,;.���Mr�C�����t#�����z�J��S�����JlP ��ʆ/,~ &���b� ��?W��b���$H�dwo�:�o|�\��ӓ255%�|��|H�v����nZ�[Lr�,��R�᐀�*`��l�\����.>�)�,k�g�&E��ư�~��~nZOǽX�ލA�P�Y�>LoԌ��i�`@�F�=�t6%sK3���,'�9)���+��Y���)7�7(;A�Lsx�C�f�r��*�X�^</�����^ow_��&��LE$�(陮TX������'N��Ĕ���Q��ggg_��v�ש3�����l���(����&�
$��\*J.�a�N��HQ=#>�쫶�8j�5*8z�Fx��h� �3�ü]y #Z���:F^s̩�'r2;_���)�?4'����Çek�*�^L�����I���U^��[��ϱ���%����u3�HJ���H&�j)y��L��裏ʡ�C��#SCT�Qg1���YUCjU�CMF��lNJx>p����r��y�u�2������M�.e���{�p#IQw��n
(`�B謉��熓+o_��.4��⟿������P���o�I�U�a)6���j���v��+�C�@8��K�P�N<�.�� ��^�zy��� K�'$��Pw���|�*72x��JI���� "k�[�lj���2	�
g
R,���aY\9,�X W�ݐK�.��榴���2?;#��	������S�z��H�ULk�sK|o�Ce|gs[^y�%ٸySF���Xt<�`�Bj*��<�����BA��T��٥1Պ��L��	!=rhμ���Z@��aDם������~D|�1����n,.�/\�*r�$�cs��eyy��DV��A��ڿ��5�rPGź�k^*y}�f�s��#����GV�w�`�a�Q� mw)��������FY>��������4�WΟ��/�ͫ��MB|�����Q'�;    IDAT���;p�,e�`�%���ǧ$M"�x+�]�,��A|F9�>�ҥ�бeY:� �����{���܌\�rS�kMI��l�h�!����C+���ü�v�5Rl����ޞ����"�AQ\0��$��:�&ea�L�'��ȅ@55>S�fx}���(AX>;]�L2��4h�����&^:/����%�՚�a���]� ���j�F��X�

 d2��T����p Z@��z�軏�<����ww�\����~�o��`�����ʰY�~ 	?��l@ubj��i]T<yຓ+S
Ќ��1�����<��'��ǩ)%㲱�+�^��T��5V*������J�!�2�63;'��������hl�����Ɔ\�rU��nJ�Y�b!�S����x3��\�٪k�FK�!�?�xl �����l��7�������e�jK
���r�D�pn�Y`PY�T��j}���f�f�'&"rQ�V�[��-gaƎ_j�8�g�	{8�\�@�����+gzHN�>+���ؒ�7o� !8�K$�S8��\^._�,�;�fӕ��ZU�6�h�J0,�T� ��a��O���,�i�:tMj4Q��H.�B>#�BQ�î�lo˭[7Hy�...�~eSY��L�leJ�wv���������5��Ac�p��J����b�����VEX��"}! ��叽��S�=�9��6*鉡$�I)L����#r��ge��1�)y��U9��	���H��mjjZ�9"��ŗ/�����n�n�$q;tR<�q��١�4�S�X�x2#��x�V|���l@�#�N�,�'�f�tI���i1���L��������˗e��u���%MM0��LW�ph'��C^b-������%ɔ'�S�G�y��}?����]o{����@���8�nK�^�c4������:BVg���@����Ĥ4%!�aL����5o|J����o��V��/�r^n�mP����S�MiA���NG��^�)�4Ha ��2� �F����ٖ��7���-Y�٪��:Q*���T�&)�����~l�RU�c�M:��Ak܀���7������pp���%$�� ]G������	���������C�7�!�:�B�iw��t*��6&Q#��QtFO�YY=uZ�}����Ge��qJM���������p�V�3�m��K�27]��&x�`��n��<9��^(��"8�{D��VS�v�'պ��m����4�U)�323=)��s�N'X�q㚬��Qނ{�Md(њ��H*�+/ /��
;�P���4@t`��b�P�H�j ���醝�R����h$��i����#Ի��4PMO'%ȥenyV��Z��yHN�=-S�s�$�x��4[}΄o4�:BZV�YuF����������Ա���#��r�<�P��X��
h����EԀ]g0`�����z�{ean^&�*�B�\�����F#AR�2� X^�t���ڕ+�>�J�ڐA��2�a�$�=�n�k@�1�>�ۙ��&K�5�Z9��++����g�.��xǏ\����;��-vפ[;�\l�Au��չ�"�y�B+p�tss%�-J�AF���?!�>���''b���/]��_xI��QL�d�N� M����ٙYY��nQrh���4M���3Tⴣo�\H�P�q���r��=lD,�\.C�ύ�i(@�����z�H��Q� w��|M�]x��# 2�N��D���c��f�@�ӳ��Ԟ!5�K����ٳ�9h?��"#����.�0�f�R��#�'G2�%_.��=���G��~va���s�.��A� �E�tϑ��fՌDJ�����׮]#�s\Y"u�)�дC�Y����D��n��� ߘ�����R�ȱ��~KeV�:_ R���N�TZf�g�E�|�%y���ɭ�7��l3��; Hb��)f4���Z>+(��l؝d*�;�HH�x���IiP}��GF="'Μ�{�G��L[p-� ��H��Fj#��C�2�E��>��s�֡��(뵝���	���,x��dJ����d�}���[M�� #
M1v��Tʼ��7���ZQ���2<�g�����x����ζ�ַ	��!�3F��	��&����y0=I�9�%�Vfz�K�~c��}��ַ��ݻ�H�O�Ώo���w�n.��nHso[��S���T����e��d�f���p�I�0�C�9I����O��,;.�<��jؕ�^x��9�xDL#;M��h�R�3g�ȡC��=ꉯ��=l8�j�7�|(�ǆ�F�}��U.�LZ�JK�MF  �#+@�-�A��F�T&�� ��7��o?��z=�I'bR����^WFCL�C��t�[�bæ���S9I�s��o��G/��wsD�4�gX�9�t��7�P��Χ�T�������BVO�a�����r��eV8uv�P�{��!J=�bxE�P��0?� G���T��WՖ�V�z�a���P�O�=%.^xEv��%�	�/��NI:�b5!d���&��u�;r��?��r^�����示��j��i�^��ڤ��U��ͪ���<(
�ろ9"Y�:T��gѠ0Y}>#�b^��:!�>�rbjR�ͦ��܇�m�4@	�B�p߁�<ܩp�Sٌ\�xQ67�y>
�6/�|����z8r>��6�c���Gt�"��-��ْF�.�A��7$�.����ΙNW�� �ͤȉ/��I�ӑ˯�"W_�(��n����4��%�H�8�'
78hp�Qt��j|��{j�SY>��G�<|w�B/���O���ʋ�%Ս���ui�m��(t�2�HW7dA�uJ��0�	�'%S��Hf�fe��=������i_�-76���}Cο�2���fcD�u�Pl�'�|RN�8�����9t�R��?H=�
�*v��H��-�
�K�/J�Q�R��S���,	̒���,Sw &@�4���|�Mp�:t*y .\�a*���G�|dC���ņ૏녟!��K�	�G��"6�8��[	N�0ǥ�uO:Я�G��, O��<������aJ^�tEv�j��h�!�$�!����0�\%����ϙ�N�A�wq��Q��#u9���fH��`�&�/]��.I�Ug�z��,�ͳ�
	��h:z�s�#t��G�����l�ݒs�_�o>�]�ɴ�z�]�A���O�AU�vMDj"�Q�����8ݵ��U��6�&��~�8=%�O���<o<�!o^k��^k���5�y����7Ώ�`�<��^�P�uGd��=��oN�)0��s�uj'�FqMb�����A����K.,�����qgo_Z��{J}������<�kW��Xs��il�Ik_z���:��g0��][,�i�2�.�%U�@��򙳿��S����5}<�ɏ�����s��n�ImC��]H{����O'�p���i��YV�܄Œ��I)-�����'��%Q�� !�Sݗs���+^���k��i���\��H�he��Mo�JeZ]t��Yoq���u�[-�Aj�H
@Ѩ�dskC�^��1���q�\G:�:�i�0�( Ut�M��]y����g��	 ��<�h�;ͤ%�KJ>3�lUv���i$���ـe P���pS���ٲL@w�~"���'��3첀A8#����}\�Œ��ޕ�k�=�����ݥ� P���c6����R���"Z�t��N�� +��/��=r<#E7o^����es�,�VWdei�*�˗�����ht6/��ߑÇx�_}�e�ʗ�$W/^b���RD� L7 f\evixO N|��F��կ�G�� !J $�H:~gs�|�=uRz�	9z�Y��nm�$�.��v����B����Fq����,h�2˔���Q��rv�@^6�Q�"U�J��B���`ʀ�[�+:�=N//���<�w�\�!U�X�8>ex�"�D�r"H|.�E.�t^jp��ۓ�.��]	0�:d��	�6�*��d
>	i	���S����_]<}���wpפأ��}��������U����]5H���C8�!)2�xN���C�9 HT�!�	 �M���|X��X����r�j��ޖ�x���ٔF�%�:$=:���fxxvL�M =l�3���&�A��` HX��[?�OvGl�^�M>�҅�ܰy�8���i6�F���
�&��� ܺ�.��Oʰ���A�UolN�#�rI)�29H>?�nO�*9�d,��v R;Hm�h d����1�Ul���VR0���Z	g��Խ�ɉ��Ic0���ی"[�k� �,��p.g�N��
1s�V�ry�ิxH#F�%���D�x�����yx�X�^�>��[r��V��ݮ>rH�f٥s��Z�u;�g���T(�걣25Y$_���N.�Y�����ɠpN�NJ6�Ʀl��1�Qd��qE��=��lk����h	� � ��r�}�ѓ��Ǟ��c�������ܼ�F����=��ͦKĄ�(>�p8�\ې�`(3�s,|�S���	��9�u��ԛ�{(#���$	뛦���X#�������U�<��ea~�*������ۭ)%���DI�*e9���5{��ey��d��-�no S�3:]�A�J��ݕx0��9��J3��#��t�ꣿ���w@��{>��o=��_Mwv����Xl�*`L2ŖQJ0��b�q�#Sy�MN� ���DY掬������{�g��-Dq7o���4�o����+�!Oǉb����{��c6��T8Tv���*�WC:�Tz�y�XNNzkT� �ĭ�y��y��2ٔd�4_{�\��T1<�U�vX |[mvy�����Wl��`��bubj�3� .�ɜ��d%��#wU�TSryKHu�%�ݞ�Y�����NWd������CS���#G��~��>�3Sӓ2�0�j��ٳr��Y�:�Ʌ�7Y]ET�ǓGͦ�Ih�a�D�ؐ�n�Q<���'OJefN�j��]$ �(��m����6�R��-5Q���S��K��z7�]WG��p(�AL_�(����9��<ͯ}���ܳ�JmgO��aع4ꩉ����/�bqar�����k��3��8�dbjm�נ Hd`͇3� +�'��7�Q�%_��V�&��^�[����N���t�1���R�C�/�Zn��S�X��!��������a�G�|�yؙ�EK��nKv�w�٪2��f�<��=o�쑲�t���,Bt�K��ӧef�,����3���s�P٭6�jg �<���`QדDГ ��(p���0��d��Z:u�/��;����� �(_��~���|������x����r��?7�d��E�6.�p=V��6��aw�DV2�I�'Ӓ����Iy���"GN�#� �W/���mrH�7�݄�c�������L��Yg��T�Br�D�ҏ)���N�H��IERSW��gu�?��?���29����r�$k�(҅k�"8��?w�p�����
O�: h��ꪺ�  '�)��LK�ؗBq �����E��zА~���˭��V5+�D��A��Q0��!溤������¬L�NI�T�\�{�q9hu�������lnl��,���s�G4�E�gj\�*S>��=�*��R�S��PE��mK�=��2��y}7�������UsXW�:��-���ǎ��@z�*g����ʊ,-�S��g�.�=��]���h� �TA�C^\+t�������xM�#���E��t�%^(Uh���,��u�̗��ֶ\�rM��v堦�Q�N��������S�z��"���2�\��kd;���XK*#�; 2z?�������&蔦ژ�{���z<P1���^��C���H�vG^��������C6�����'A����C����@�4<�3��$]��/�:�-�z�w�z�TL����O��>�l�/�ѿ����B�P���'řnW�>qh����/�U�DF��@����R9Hd��y�����[�n<&ϟA�\��s<LȬ)uG�w�do�@�L�)��사=&��'X���Ч� ��M��K�*
�3M4�ԍ������)��cG�w�����V1,gmw���n���j�iUҮ�)�@'"HD��|�d�BA@%�r��M��rV&ʨr#�ږvs�3��ё�[8��� ���\��s�d��{ ��d�Ȳd��ēO�ɳH�ӓs���Ǝl����A�Q�g3'8
 �M����h0�9v�8o�	�\�]��|����f�64sFK�w�y��+R��eq�����oG��@�0�m�%�s�DIV��--�x����g����7	�pJʠ�$�N�d�hC�A��� �1ڗ��O�>� ��>�T�K��C���Vy�ǥ��5y��%����ɂ�U�XVZ�YO�hgT��c�.
`K�+����q:@bȖQ��l
0�7���qO��G�H�F��R�K�Q�\&�CH����*��I!�%/�r��Kr���R��&@v�DZu�c��4C����ٔ$'�����.�8�O?���
 _|����}�}�����s���TaԔ<��H� 	�t�  ɑ��)	r�IK�>E����ʙ{�o��^^�^"./�?'��^b����*��K!b���'ؕ�e�����ʬ��猔�E�dg�^����+���j8q��.|�`bl�+���V�Eyɉ�U9�ە�ϟ7� �49O�����a���C�n\�,[7o���WǺ*�B�[ȁ�KJ*ݑJ%!K�(�������R�l��dw �6$Si!���ڈ���Uk��nܹ�9rbUr岼�Mo��#�e�ђ�76�����S��g7���)*ʻ��^Y��Tf�x�(�*�Z��h
<q=)Lf9�����ҥ�dog[���?�lT,8K���x�N��ٙ
+��yo��v��=﾿��=�>sI�J,��`X�8��`*e���b�)�0`d�U���+�b� q0��!�@�Z���]���gz����}M}��9�-L��j���gzy����<�w�}޻{�^��/��[�,��xH�"õ����пJ�"�?�����?�Rgl!�2�ǁ3ac3s��3o�o�/��]~�M�$�ޣe�}��mlm:>��ƺ�#xB%,f��R�$����/מ!M,�u�P	a���-�a�Gǃ#��*��2��>�ơH��Jԥ�V�!��5���A��}��-�~��V׬�PImϬQSo=A5������v���h=�݅�Wj���_��o���_B���� ��'��?,���\��N�u��� �v�92�v��4����Hg�`���+@����}��|��͝�^*e�-)@nnмF�݁�ܼ��y��ݷ;�,�-��Դe�9�� ��'�M7\� ّ �,<���	�24��"[_�TIݪ�49�x漵;{��W�����6��	h��V?ؗ��z��mm�d�4��'���9��T�I��J��d�FF��Մ�ױ�W��m���N[��m.*=yɉ�Gǵ.�����0���������_���\��Z��-����[$�F�T�J岝={�Ƨ&��M6+���J@60٠�*�0H����TE�^� �^o��ȥ�%`@+�XM�k�����{od�d��c#655a�bEfj�~�E{��W�w�Pꎈ]��s���=H��=�b,Ke���c9a>�I���/����E{�k�ξ��^}�Z��=XY�[��K�qwG��B*�	AĘ�r�Z1���Qai���wes@���"�T�:y�I�|�� Q�:� "��!�@٩����p�\c|�D���aH>O#<�������z���,��>���bi+ab� @°b�1<JU����=y��O^Xxۯ>������_��WE�|�S��_��?ɷ&��Ha�-k�.YcJ8�С���
��$�Q%)��g��O)@��,8���"�P��w��'uh�O=i����g?��cHCo���v����R��ӟ��w���FX.�D]�!@һd2I��A�?g�OX�ײ�7n��ֶ-/�$�^    IDAT/���Y�k�6_}�lk���ꆾ �F�U!ڊ�4��+�v�쬝89j�"�T�[v��c�VmscOx�f}`��bx�d-�)[BP� �@��Pwhs�L�glr~ξ���N��d۵��~�l��"��MĵaPC�,W*��%	(ܺu[�T��������ч�*����4�'�ڈQ��Fd�D.,=r[��-��ްE��nWV�|�K^���V�{�����1	򎏌Kjq��/���F^5d���y]a�-XT�����*�Hꌷ3��{�x�|$J�Ik�&r[8u��U������
��
��do�;�?��z�Ӥ�:3;+��~����숧焊��Jz)����Np8tJ��a����I31�%@������I<>6�������ŵ��!59:�2������q�������kh��Ab��A�P� �� �-����Ή�W~��3o��g�}��˟��Zz�3�(�>S�D ��D�H2Ȉ��_�.�	v%Kf�jZuv��>��k�۬8>a������������e&���M��ە���z�o����j{5�N��Դ]9Y%"��^��	�'�[���}F���z�2jkcS��r�`ss36?1m�^��߽'����z7P�(�Գk�lmy�ݿg+w���j(����X�<l ����!;E�i�.\X��)T��֬������+�
 �j6�k6z�w��U��!P�jH8�?�336j��^�$�8r�ձ{���m�n�����W���>��]�tɪ��v_֬�u�x���u����H���8���"�Z��'�ҡ�����fS�ls��]�x^=��w���?�q�a�!�_*m�R��)/�s�-?Du�5�{��?�S�j�'� �8���.P������e5����O�J"�� 9 dR6�����v��e�8u}�V�6ls�!Ɇ�w��P�>��	�>sF������݁�+�N��ČO�7^� ʞ�a�F���%	�*Ç=e赚�`p@SZ�;w�N�/H��;$  ]���� �����`0�r��m=X��eg׺�du�^�`}KsUZ ����K+NMn,^y��O]��_����r�W0��+� ������{�+v�'
���hB�TP�#��!�1C�	�=Q�B+�0S����v��g����,;:jݤ�%�v��k���b�B��F�699n�.���Ș����V��D�01v
���d�����>d�'����O��X�`\�N�!.,Ay|d�V��ƍ
�,8�k����]�C{�ݽon޴�u�:0��g��v���d�g�R�N���S''�TJX�`CG�ޮ�m	#�Yk��v��W�~�	zG�e�O����f&m�Ă]�v�ϟ�3�Y��v��|�;݁�%6}����#ᷟ:{F�k��?�������<d�J6�~'���2u��H2,��<f6wvmk{[:6�Ϟ�'�^V���O~�^~����G&��=��
R[��O훯^W��	�VR�=r�>�B����!��31�T�9t�0�һ�h��B�zɄM!������ /]�!̣��mm�*@���(�L���P���z��	Up�~泟Z����Ą���Ʊ�e���`��'�ۇ�#N�h�A�0(h��g��d��~׮]�f��
��ۛ��V����4`e��1����kKK��p����`k���}�3z�D됍'zF��u�:j��镳�����gO���k�p��_��WA�&~�?�}���g;;��������9KY�('gC�B�n,j6t�d�D�R�K�6GP{�iH�ؾ��N֭X���ȨM��������-؟~�9etL>G��L���֕>YL��sd��$1`�(OZݎ�a�H�!c��ZPEQ�"�t��i���;(h���u���~��22��9B
P߰Ҽ��S�b��8���@1O�HpX&;������U�T� �c��!* �6��@�}�u{�<صJy���"v�j�ݓ���͟�����܂]{�[��Oڍ;�,L��u�b��Ë��Tc(ei[P��s���5�up�O]{�ʥB{ ��g0�/�À3'����mn������F���T�����Ο9+�(�/~�v��=kt6::"�6�����M�O�$|�/��d^�X�FQoU�����ݑ�!��?E0p�pO ��=M珩���I-[-��̬]y�-�u��Mv鉧Q�m�mG̓}`��
�@K��
���v��Y��7o�͛7�*�*Z��z5�=��V�ח�)�HH����`r�t�k$9����h����Ta��Z_^}d��ܶ��M�iq�K�K&䟽r�����Ɔնw�Z5K�[�'����[���ء,R�媍͟zp��ww�g?��w����+%�*���?��/��ٶ۾�I��c2��VXAZ@W�E
VCtS9�&�-���삝����o�V+NM[?���6<�G�$�6�$�E	��Cel�&���K/�����jy��霘 �r6���M��AIE�8
T�]���BIGI��+C��(#/�;/�3�}��/!���:}����`���`�����W�>���˒��˲�A0����x�&&�V�$-�CҞ��h]-D�!q��C��e���l�TI��`�q�7|�\F��S�3v��Y�N�ړ�~�u�y�s�Z�.���mo;Nϙ1	�¯.dU�ݺ}S"�d�l��Ș�H�3\�v��( ��(3�@E���r���ml*����7"�dL˫+���۝����}1>2���k]F9�?�W^z�ܺ-Q��^M
AY�W��Up$�V����}��[m� �iq�)�R5b��?a��@�4k���!sf�.?��=�_o��~�RŲm��m���6w��� ɡK���<@N�L�����
f�߸�������ǹO�
׀���a�~�MEP���D�� m �).����.���wI�=����ֺde�����kY��5[����5��S�D�nI2Hc�9�4Z��ߢ��PR9�p����O��w��������llԣUȏ}�~߭/~�Ù��d	>q���Z\��"�$�l�f��ֵ���V��lu��_���g��M�=� ��wm}k�^|�E�)�i��UF�wds���*y,V!����hJ���+��c
�
�2��G��d�Hh��l��d�AS�g��["�3�Y����p� ��k��/JIGY�#@ܝ�-[���.� � ���)��]eF�I:��ͮ��L�+p�Ӗ/��Xu�	�R�C��BY�m}u`�]_�^�\�R� :'C�b��J��f&����V���g����j��]��?P��<��0���h���(�r/��gK��35;'��y���k���,�aG���@��=���Uq��!0��Hy}��Y���j�P�ӗ�s����W+��®o"8 &���M{t���5z�y, ��b�Y���5^�*N���z ����'��-�S�aٔ�ONKN��'��Vy^o7k���-+a��W�tX?� a��Qy?�h��3�r��
�T(D�%]gY���M;c�	^�G�Θ���٠ﹹ��H���Lv	�&}�b!��@Þ��nܹ-O�t6��vP6��a�k;���~����?;�mڰ]��+4F��#@j d~t
�͓���o�����_B\<|��� �+������������#ɶ;��ue=��A5D��O?��>S2��
��҈��,Z�T���g��o��O>e�\ֺ����v�K/��f2���^�h}���Zmo�c���kA�@M�L/�M�#aב��a3p��Z�)lbNO�E��`c���	;uꄰ�mM��v��]�C�jJ���t��u&��ՇK�CP�z��)�zc���@�%���W�����V)o[&7�ɉ���OK�b����A��3v���"���R"�*%��̪�#�x���홯�F�L��N�#��ɩ)�o�y�,WW b	UP2я�����$�7Eֆ�������S�*S~��O������Я��({l2��۽��'gT��U�,�J[�Ӗ�
ڈK�j�Cє�;fS�C�궶�a�޷��Ug,5Pp�Hpn��T"�����!�8� <۹����I�e�!˄x0L��c�����3g��Ӯ�4w�5�={H`�{��հ�'�ד� �Y����kw�޳��u]cd)��#h�6T,�ia=�^�v4�b�����=Jpĩ��������gm|dT=&<���ݼ}K_� �\��A��{5�]Y��G�V�\���Gݬ۴L�4�2~��!�2��@2�����M,���x���������*�� �S��k���GS����T�=�-�Լ7�(@2�h��(.�\tW��O��M/X�2fc'l��%���g,?Z�a>c�V�^����q�u���Q)W�(��&�V\V�)堦r���q\�K
)y�G�� HfH�6��~&e6����zJ���Z�^y����>j�L�;��m����;�le��q]$�Ȟ������$	�}	sG0J*�B� I&�͐}u�Z���4�Ͳ�w�D�n��~����w�3�.H�`��q!�Iyy�b'Ο���i�����̂5�}���,�6�gk�1�d$l�TM�j%�u���_�cْ}	Y����>�ꨲ;��t�uDp��14ÿ���[a�Ӱ*���� �$�'����_x�[�\�0��"@b����#�\]������ؠ�1�����F8�<�#�)�|���a1+#h�?�9��z���j����#657k�/^�'�����|Ւ��=�XS_��j���0C��\�|+���bwG��m���p���+�#Q��댁C>j�ɡ-T����������o�R>��.�ߺ{�Kl��ق�gЉd�M�����{�/�uۖΆ` �Ǣii�i�}%�τ y����K��[���� ?�џ�o_���ϙ���H	������^ؘ(��������9��a*g��)+ML
�327oW��f��NIQ�e]{��dϿ��i��JŲ��������꺸�H�n��A9}�-�p�NS��awx.�h#S*X�ӷA�ҫ��w��9�ipS���[^[�7n�qp5�8|  66��~MÙ����U�lV�3)zs�9i����!+�u�A��&$Z�BJ�hV*f4������:���v`��VP *��e���m�a�H�4R�gO���E�?{�&�l��ۃ�5��!����k�k�Jz��/�JY=A���Ғ��T�(��Ⱥ�8�m2#60n���(��WX[>��@�������ܹsR1"�e����KS����IY�����hC=���kQ���}�}���=��(zG� uxj)2fd�/�4HM�� sUC	s+6:5a�'N٥'�ٹ'�������l��� �d�Rթ7�#~��A)����栢�!�E[׈��vQ���D[���e�i5So�������$S��.�?oW.]�|��d����ml؃�{���+1(z��j���?[k{�;[֩�u��8[z�4Nyu�9#N�A:i�l���6�p��̙?�]��#���� ��??�S���/}򗲝��4iD�E������9�:ְ�y
��wer�"㛘���&&�̵'l|a�&�fͲ)�o����=�`We'��Q*�4��]J���% #�v<W��f]L�(�"x����,
�1n��I���ĭv����[wle}C�	�-�W�{g6���֎���K�)�!@R�9$�i��|�cX8F�,0`m�?�Z��RZ�R)80��V�k�[-�ucIYy����4N�LƁ��(��f���!��R�L�N�a[�[m�zC�Dt�cCI\u~F��^zU_��H́��ʒ��d�T`�CL��������U��X.��D�d��5�����{���tg�~�� 	�O��Ξ��X}{��0�j�Z��I�WȀsզ���jCb�P:KE��EU �w��B?w���1@j�
V���9;y�]y�����V�w���;R�g��H���:�k�`
.
°Per��{BUsH#��pAr�B�!k��9�32���K��UÀz��U7�K��C���]�@=���k�=�����m}Kï���k�֡��BC.�h�}��,Q�C+� �d=������s�����^����8�=���̗���p8L��/}�{�^z����LkWSl�Y�&
�5�9A���i�ű]�"��9�LLZY��1[�p�&fmlnβ���O}�����WJ�r�v.o��J��K/�,��F�)�7^�,B��+E  K:����٩��R��a q���� ���myuC���`:�̒��w�k;M��XWp�>���rKJ} �����N������a8��h*�*)`%�'�6:Z�� ɠ�Y�K/^��$6:�*X�R��s)�������r;u��,��� a+�;�o��lZ	i�l���G�����X.������W^�^��<U�ݞ5�m|S	�� ���Z5}�6�p�~$�����g�-o~�]:{Q��p�N3�(-
��:mv�E��;���mXc���5k�k�k���66	��C�_��1R.� MЌ���TPǉ����ę�!�	���X��zZ��q	�^{�e��q{��N�3�f�]
��9�1����c��k��|*�(��*���vxJ<C?8Q�X���'�^�'�^S{$��԰o�����z��H	�v����l����[��q6lXb�3��--f�=�Ef�M)@��Q��Yuz������<����o��#t�W&.>�WG�����[_���inN��O�*z�d�ꂹ�_v.�d�;#y�[�߷\y�قU��Ub�#6s���/�[ilD���%���Q��VFt*�8�p¦��-�����������@2RK�T�P>dF �[)+#a�n���=.��ۙ��XRɔ՛-��]���n�˺�=�^�e�f]�{[[����<@9���Nd3�".��$K2�� �V6ֳl }K's�H�� l"83�VUf߻�l�&P��Hb�2��K��¢��L��Ԭ�'&lzn��O��n�K�A�դ����);:`!�~�K/��/�j�RA*04S�6"�FeaC̺�
*I����C'Jiq���7م�筜/��٨�V��ރ���w��^�.����y����5�U�[�6(j>�I���C�	�ǭg
�&����b�q�D�h �u�{�����͆w�=yYϜX�����;w�{��3D���AՒ��.%���z=���U@� 	���j����{��?���MJL�����A^30�s�ϩ��0�,ȯ�Ѵ��}���QX��ӕ;��Sk��ښp���}�9���-�n�_)5h��k��#@�P�3�2t �EKUF	�K��|�Ե��<���w��_��WE���_����>�����d�w`�D�R
������"�g����*�Gl��Y~���d�'m�ļ��G�+���n{��0c�9p�+e3�72���py�����n�d��EW��ML�S)���RH��m��lA���,e&f\Lz��_Y[��]�X(�@�logW��e��ZM���e���h���:X߲)
C'�9+�/|ې)a�,�MX:�]�O�E� K�>��Hp"a�Oft�5�٤��K�Uɞ�*��s�%�e�ᵒA�W(	4�R�MWo�����ޛLelgg�^���3�::��jʎ0����lf��>�����]l陓glvf����F��!��2�ߍU�?,c��P�خխy�o��=k�X���l�V���0|B�Ѐ'�Ԕ�
�a�{�l��Y(G�*��f׃��,Ii�s"�,����%����'l|v��N����Iy�l��x�"�&AX�<}JZ��YY]�%r�$�E�3�^�!k\}l���}| �'��_�p�N,����zA�b{�@��x����z�qPS���<�zÆM������Aa��G>JII�	:���	y�Ab�R���?w���'��w�_���w����g�[�~�2�4Æi�k�M�ҝ�R��Ƭ�NZ�ݱl�j�Tֆ#e�    IDAT0��-'zҤM-�)��bS0E��V������LL
~��w���e��'������,-�-/K�痰b��I7���E�ޭ��(��''��{��&�e\�X\���O}��H��`oW���I���:��zɩ>�����L�]� )vv�}`����2	�fh�9�\�AH.��o���5k6�,�����$W�EO(%b2�rQײ:>a��361R��|�l��6?�(�(�SNp��s��y�t�nߵ[wo���-\�|�*M��kUj�b&H	}\hmd���Aw؟-h�Ð�@���H ,@ӿ�z����a�P��ޗ�5_	�Fd�ٲ!�h�I�)XxIM�ic�I�&nd�1�į�c6	�O���`�NO�'�X���[�.c6g�jE�s��̌�d�Tk�m,���M���c?��7��u2����o�Սp�����u Uơ�=���L���`��/ڙ3�D0�Q�����!r���hd��n����mn���Dq{͆[MK��6l�,�\��l�ї�j�/�0� �9����(4⻳箾��s���d�W��O���/>�����D� 9t&�c�����4�	(� �雂]2���dE�ծ�,;2b��qˏ��)ndj���3����|�l�꨼IN�̉~��lг��g>�Y_P��zg���|^�#�X!,0#�za�U�e;�;���a��d�
,��eQ��}��{�������$��6@9�2��N44�� .'p�
\���1qD(6Z68p5���D-B���-�9�V�P,[�3���u�כ��e���u�e��*U+�T\@ 3����ϝ�*��y�<acSRPM�5\[[��)A8�xolo��ʲ����!���ɂ���j�\����MF� ��3gE]T���(oM�$�G�t]k#�`�/���'Pք)��mw��^z�d�	)u0�uRB��� UC�hh�Ș!� �v\XWx���'0R9����E��uz�F''�0>�L�����[-e�c�=�<i�/\�ΰ#"�6b���j
��5p��?�k�- =��7�P�'�V.�yW�/+�_MO�+0F瀗�g��ە*?C/z� ��0ba��ݵd�c�(I�a�n�d.;D��#�,$脈�U�]�(]�ѹ�/_z�������q�b'������ҟ�\��RCj���Q�R����'���C���&e�%M�;ä���VG,]*��LMZeb��dp��#6:6�qnj�h-�E�F��K_����Ǳ8:A��#L"%��4*=Ͷݺq[Y�@���L�0?�e���'+�æ�@�hgm����p��W�j�F�R��}�J`�Ė`n�=��� �Հϛ�;XYi5l�EWF\��l��P�UKU+V*V.�m}s�v��*�)C�L�����)�P)����R�
�v��9{��Ӷx�]�9�-��澸�`� �z5��b��xW� ���駟�'�=�,�罝�$�k���m�4��P'� )��	�<>@n$ck��{��>��kx�NF��ɴ�҃tv��3x�d�4Փd�%4
�T�%0)C�p�(����@�$�%5�����u��Gs��;ϔ��^<{V}`z��jBA�d(�t�ϱ긄P:����~���t{�C���2���g�ʨ��X�P���R��Z,UT%�ˣ�;z���f��A�݃���8�9�t����ή%*��
���+���Ӏ�X�$���#�+Xnl���O�:q��{���� �+��3������d�q�
 �؀. � �4!@v��g�AerR��Lޒ8�14�D����䴍�&flzf�&��l���Fm�z�^}�����k������ �Z����xX,n�T	x��iM��߹'5�KE5�;�����oޱvቔh\�}��`��=mZ��8�6P�DfKr�"�9�Z��>�C��Y����GJ��6c������?�� %�&ɲ9�_2*;�.���+����;�=��[���V$�G���������[z`�9�����ݖ �;{�Y�Moz���dF7^�<\�t����!���#��}̬���넾X���͆�b�a÷��Q~w{
�I�t=��셃�ѵ@ݨK����� 1�>�7F�L�� Ct�Z�ih}�7e���xn��F��*'�P��<Z���ye���x�=2�n�OHVn~aQ�;d6j�h�� �w�$gx��Xcx� �8y��2��+��Ç�$�!�le������^�m��b�S�,���E�6��k�n��ZuK�� ��A-#�O8�P�����(a}~�0����������o�� ������;/|�� =@��`.ua`҄��⮄11�``�DI��Y&kd��b�@�D�3"~��ܼ���ۉ�gm>i{ow����ko�n��&L�i�钔��=��G�����2M�os����]��ށ����Ɩ�S�bV=��9A.n�v�v�8U���Za}�&�nG>��(ِlR9���@�á� �	��#�&�]�TZp�#��\v!�t
aW�}�2���iwo/(��P�g�.@A����Ȧ$�@3�!@Ο>c�/]������ܼ$�L��r�������� � ��*::�)�)Ҷ����5���$�ē
�H�=\^��-�xރ������R�I����֯7m�ej����8�G٣�	��#�'���8,�ÚhH�Kjck8�:�\�R�h��9�^2!�
�
���L�1���T�`_��!��مEI�gD"N�=�CN��@��}����H��\���z���d���	'�֩�
W�l�7�"�	���V�'ong8u%��5g �!�|�@Q��tkWd�����ơ��m�?��2��L������������.�﻾����/ax}��Sl^ɯ���|��/��?�vv'
�K��B ����������3!UeJ:�B�D��oS����e,�iQ:+�di|��g�lv�>sN'��ؘ�l���m��2�c34;><PI��L���/恕Q�Y��ƽp���|����*#b2	�ejz�v�v���l��#k7;:e�l�7�w�U�t;�i���YT,���?(�$�ß�(/a��;z�Hp|� �$��ۻ�Q��������A��a7.���Ty�T.�- y�`��q�LL�n�����:jа"M�H�F������*5;]+`}�y�H�kI ���Q�;��/����N��H,�K؎޸uS^��V���^f�QW��^��Ы[%u�<"	�0�d��Fկ��\K�/�#ט )=ȁOڣ�y,�E5����j�!�ۇ7]Z�����i��e����3
��RQY;�N�cTCH�U��d�A�Y9)�Y;�|p�:D�������Ǐ��)�����)�&����" B�N>���N�&[���>9<� S�
������m�w�ֱ׶|r`%�G�f=�>��@b���O���$9a ��0:ac�^[<�=������ ���w���O�b�ט*Y݆����O#<��~ �sb��NY�!0/Mnc�@�9}�LR�z��e�65�hgΞ�9A)fUS�� �t�lnNG�dY�+��9�2��Mr�K��B�Qف����X/WR�ܾq��޺m�}gmt���zeP��g�#e��{�MЎ�1gR$@�SQt�]e	lZ�8�s�!��h�>H�Җ�"�)�D<"�d�`��=�%�/X6�)e,?:!K�r�z�'�Y�W���I�����7�����E�(w��a62��N�Q��Ct����씲u���7d5@`$�5���@�:d���^f�*3lw�j0i������a�Ll=f�܃��|��Mv�\eZ!����21\w��A�!{�kU��$+�EH���%��§�jӰ~�$�f��NN�Y8�o~ڦ��,�Uo>ln}͢�����xQeaa1-'�E>Nå��re�����ف`F�����5��׺�����p��.-�M>�L��M��W`�w���' �TqM��p���v�IP��F�(�m���_�?w�=o���c �~����/��S�������Z�br��� �Z.|���&@r�X|"��i̱�ɛ��)�e^��L�*SvJޑ�)�u����M�f�gr>Y��h��ͦ-�
�9'(A���G&�de�1�i�ַJ��j�t�=�{O�f�f��`�PN'L"(��1�� 첈��\$r��T:R�f�C�Qߐ!ST�3���C��Bx=e3�?�>�J�H���P�Ye\�1���5pe�#
�8�e�N�+�I�H���X/�+R]�2#�,��F:�z���'�R�Ix))㯭M����ϟ�k}���3�*H���������V�'�U�7�H�A�� �l1P����{�{A������S@ψjǲ2/��V���)�{�C�w�����-�����}�1�B�RŜeJe+�Umz~�N�=g�'O[�\�`���P�l�U��B@6a��@���5��|�(2�RutĒ��z�(�c���8���4���hh-�c�1�nv�S�K@D�l���B#�re4���JL.)��K��g+
f�(zkef��⹫������ǫĆ�����_���?����S�ή��a��$��,:��JD�)8b慕&.m��d�`��%K�9�Tǭ0R�<UD1m͎��PW�dTy�Պ'Ct����lr��H*S��c�2ټp{���smom�?���"�#=���%'�A
`&��b&3ul+@Ʋ��O@s�iI�1MT=��FU �)j�C}��%�V @��ג���4�RHA� ��S>_,���'�c���P:�dJ��T��$ٴ&��
$
_n�+ss6:6fy�H�lymE�
�	��ׯ�!˄hnݶ� ���@�e1@T��CI�ej�3@aɬ��Te @~�+�=� �����*�?��[£�z�1@J��ҏ�iC������A�P?��7?C���J�
#A�Ʀ�m|z��'�ltb\��my/��}��'SW�&L�9ܵNSy�I����Ke�=t(a"��u]N����l�)	 �".�탺_�.д���8E�� \X^H�=ex�ƀHR�������-���S����x���;��?V$���_?�}o|�S�,�ؙ�wQT����A�;e�Pn�M�6�bd!��*�)�=���R�"�)���d塒���P�Z����6f�g�MH�T�H�ͩ��`\�&���'�,8,!���z�����z��{*��?*�!(���˂q�,��쯡u�� L�G��GnpC/��q�3hs^
GeL��A�2%�l=3r[ I!;W/�'�>�G��N���S��L�kN����&��Ց1������i׺��:M.��! �驑��ł�9Z�v��W�q1����U]�5[[y��ځ0y=Q8)�|�k�;6)��pˁ�d2bI������Qz������6����c�+J�q� �C�ux�^��0�|i��H�Y�W��V*:x(���s�� A�!��҃��@3�ؒQ5�����!J|ll��ƸO.����@���+�5�ܥ���v�uoeġ"A��L�]���û#��0��\l���3Ie���	+M��9q�ʻ���?���[�L��G�]�}�O~!�ܛ(j�4�=ѠG��	u������h���R�N��d��E=�(#Eɍ$SZ� �$�n��l�pV�b�ZL')(�X E���� bpS�}~#\��\�YS�ɇ���1�{�7�j��}��J���b�@���v,�����#�F�VeS�9�dJG�'DI6m`�Y)�x��K�i[�@�ů��+8�`31g��`E2�Q�L)�ϸ~�\��61埜��,�c-�c��*C���Ӫ ����Q_wd|L�44٤H��گ�|�n����>z�0)�+z�n���0)�qw��k�z���D�)�~M�WZ�V�����߁]��P[#�@$�d�����/�e�[��1Z"Уԁ�Ff�i�Y؁`e�uH�b�b�r(��+x�ck��hYH;�<|j�G���Ș�N�	�Z�V�,�j�z�w��栗K&�k�\��������\�
Y9�Y��&!�/
0I{�۱�.Cn� �� ]ͧ45so�ܕw׻~��� �����^}�O~!�>��&�����H;ar�d�+)�E����w��^�l�Ev�� ��j�%y�Ity|����"��2���{��lf�QzjH-���eںgQ��uZ]Q����%@1$�y?��JO�X�<�+Y�=�$��ǳ���AŜ�9:���>�~�a����b���HI�oڐ�׉�+� I��*�C4�OQfgҚV�`<d\�ݤ ��� �j<G���Y��.b�x����L.�L�rl̊���fzvFח�AR�僚��_����&�x��=��?�z�١�a��+��
��;���B)����ẅaN�}2hR&/o��G����������Fd)�4A�
�
�6��WF
���.�j"H�l�d��%����emBJ�	S�[*�!�%֢��i��U��u"���a[�1���ގ�H�	���p�y����2�<kd-k�B@�J.#��k,H��X�}�	d�E��Z�����ŋ���]�����c��ƿ�����O�Bi�'@;5�*.Y/�m-�����s��@J"DI^� 	��)��q�] �!�'�R��i0/B7�TP�$�a���G�`I��7��l5�L����0 &��Y�-I@"((��a�pwL=���=���~/5R�XhAUFY*���%��!�{�oboͳG�s�~�b'X��IHf��`ɆB V������5�w�y=�ac5
J7�4�M'�:D����,���{���.\\V���g�⃳��J́m���	�I�� �g]g@s臅�6�c��lYP��!�)�>��p����hE�^ [�`�T�N%}�g?�|Q�L�LM�����l��3�;�P�s��E ~VW.o�\Y_5T$ �EoS����j�bS��O>�.za.��y3����a�σ};8�뚲/ayL3�p}/���e�ҏ�����?@�R�����t�i�|�l�r� ����k���w}�w�2���|����j�� 9h�H� �q`Ɔ� �oߘ,0{5�=@j��׌�Eu�fK+�KC7�> (����S^�`APRK����*Z�����P�� �LC��㸾�Q���CX�(�5h���=0�L�L�@Y p9�����&����ȮU�j��T���gKޓ�2mC2&sI�D�E]u�CNT�k8�Q� ��B�BG�XY���\L"%&|��sd6j� 
d<E�C68���y�����T@��d���X�-�r
a��zX��v:�S�Y����K"� C��JQo�w�(z��oW�-ٵA8�|Ƞ�1�����(�8���)�`�����"�����@�0VR�U[4�P�"�{�㰅�q�@<[NJyJW���}��a�0e��j�Ym֨��Ok��I2k��2�⹸��-�0��Q��Wꢡc(���"t���A '$��d�EK0��\Z���{�����<^���3������|��<��z5vk�N:�^vȝ!X]������H�pA��q�d�*��١$�ᐪ'Ģwa�~��ӗE��	����/�)���T`Ѕ�8��7�+4�"bCGX��2�_Ї k�q��q(�6%�mеL0���%hP��g�&�3;B�2i(��T7n(/c/��7.J���9/(Ė��%)��T�?8bӌ�?
d�lLM���r�5ʊ�>� lA�4.F���78|OP�����v���;�U��^��Éo�M�^�N������)��1@�~���ҳ���2�3�^lsH��x�� ǁ���^�����/�I��4;d�v{PU?���hP��C�#4<���k�c��p֗_c�w��McKB9�P5    IDATW���J���#�7��v6Q�J�;�n)p39N�� Hă�`��բ��y�$�2�*�A��+к���Z	l�u�Y���4g�j�����'��_��O��c o޼��Կ�����?��j�3��(@�"�{6$L�>_iZ�qef����HJl6�#HM\�PdN`�S�c�0 ��� X�tҰ��Z�9��(d�q���z�]�DX�G�<"@�R�k<��
�@�Ș4�����@����U�����Tj�Vc��Ɏ(���菤���[�GÒ.A]0��K{�CCL�Pbk���-�Rz#X��<S#���c�l�Y*Q�AC0y�0|�����_�JʠȲ���!+we��Y{��>�YjH@�axpx8@�h�jG$C�(ε���G6��P&x� ����������!�{�!�(�xP�`��������^�e�!s<�hq�	����M �'��W�Uך�W��Y�z��ѝ4�/{l�8N~(gN�S�P'����7�$�=��.R<z���@Yx	�=��990�G�0�U�@Vph�bF�<dad����}�2ȥ�+��'~��K_�*�v5ץ�T��* ���$�2��.[G<%� ��� ���}�ȉ�SA�\�w�>�C4]b�z<�W�
l�S��f���i����Q��@m-.�jS@+B�G9�r�X��x��j� ���:!��?F��k
�h=�he!� �l&NaàA1M�߻̮�bɬ�.�^����1@���!�=���*%���u������:$�þ�eO@II�`?"b�
C
:pSa4�l�n��se��lr]�V8���ClT�;,h��H�?S�3�ZrdtXU,����y�x�J�� ���O�L�e�8G�a��H��I	ă���I��4$��ż��q��k�{�.3G��C��xK ��~P�a�c�ms@�E!�IB�
�e�\U9?�aM�]��[�s�2H��b���(�H��鑊�+�w�/_}����}��� W_|������>����d�J��o�~Ӓ�?Lɇ������B��)��Ѓd2H �^<�"��j����;t=Ez�*�$�5p��n�2���@����K����]5%H1���ݍPG8y*�]�y��c8㢱�����}����X=�;�:����g$���2���LB&H�:@e�g�㳬��ծ~5�^����qB�]h� ��k&dI���'�f����
�lL����H9�cN}���LK���\6�#
=���������/��{�mJC&��aq`p	�*(�
��Ӑ,�r�u�E�3�BA2���I 0�,��d�Py��z���&l�S�!PxO��t}�pe�k��3)�7�س[_�\� ue�.���K>���s3L���B�8 _�k��.�n�!��c���DAS}J��O1@��#���Ȩs�#�/\�����<^T�W_�D�S��o?���+?Z4�9�%~��Tj����u�
�b���'�Ч��J?j�x�[�bP;�7 ^m�f-&rj��z��GF���JƐ����*u|!D�c�<���AA����*��Y���)[�?)� �F/�X��0R}�E�[?P�d3B��P�5�h�P��!`cDV��K�^j(�؃N2&������}��ȁ�*��)��=�V<sW_1�+A #���<����Љ���?�&Ȟy����a�^g�1���I�I���P�����Kne���B$��x���=V��5�1���u���l� �&��)����z�:��:���5A����;���B��AaF��i��C6"[�p�+1�Mh��JG��� ��pW�W2�CT��Y@r���bJ:�p{�.�!�G휁T�T���Ӓ��#~=>ys�~쨆�O�w?��ƫ?Z�7*� �ö�Hn�M�:�b� '9|�6�� �^>6�v�rM/	t�C樌"���'���1���Ay����>Q����&�̏z�DWV���c�� T�8if�E��Q��u���w(�R@��o�=Em
�ʡ�D�:F#���W�3�P����"n6[��O6���`��B�B��r���x��un]���+��q�|��F������O��@W �Aş�k&4��x����S0Cf*�!z���E�u�^-K�l��(L�	�*��(��ܪ �Ch�/�b��Shi�F�e�ES4W�kN�Lpԡ�\��:�����c��l��)��צ�P=I��{$v�����X|�/Ѷ8f6�	��X��J���V�*D���V6j��C��\��L��$����(�"x�A�3��Le.�O��x����������_���˝ ��7���n^��b�Q&��Y��]T`(��eH9� ��F�OF�.�z(Hϡ�3����"U�,,��L��PH9�)0������rd���*�**�x;`ۇI�`\��=�CK46�OÛ� ��E��~�h��RhmNf�}��M�]\���2��N��l<8�9��2&�}x�d�ދu��C		�D,|\��T�h+l����0pRi�t7d����D%��SN�z���X=l�W�S�����*�
� �k�b�>�R�9f4\�0N� �g�eJaW�!s&�?���1%%��1L�/���C�+�l��.0���!L(wc�4�=�t��I����{p��������O8^��M�Pǿ#����`p|�0�Q�uA}��#�mDYH�ފr��|���ȥ$w��sir�K����ۿ����J���W �A����?~d��k?V���d�ؾҀ���08�^�:ÀOa��R�
��#E��w�D�@���f�ytL�c���"R��\�;��
�����Պ� �9kX��Y��0���)Xx���#�C������ �1����]ޒ>A�'۪��{!��[�&�!S�FR0� �\NAd��A�$��nuP��~���%�&���DѷR���_�\X9y/����r����nm��+��;��WVX-�?�Իd���*@�=k��˽q�41����Q��>aǇ���0!��\�#Z\qۙ6���x�(���U`
��7��4�s������]��� <����`����vܹ���:�M�/�8�%r8�BP�P,0t<�����|��Т`(�u���X�����p�xb����CK�/�i;b�!FN����pK�*�TC�2(�㱄�)�G%����r)-M�|a����}�;����*@�A��_��ݹ�ʏf;��b�ei��e��5͎�� ���p�k���C�^�2x���y6IiM���',?:f.^��O=e��1�k�7낧��:�GLW�hH��%��7�rPj�!z��o��d���i[k����.����"�v�ZuL��3�)7��Ay�2N	�d"]-�t�[�j���@!��Ҕ�$:�x�A~,�W��C�I�������~.�UtCih]�G����D�L�h��r�l/�f6c��2%���o�;��U<q{bK����Q>��]�ְ���oy��xm\�v�ҳ���=�
}/ �Z�y)hC����ʌ�8�j!�����U������Z)Pt�`VO6z�pX��(�c�R/Ǖ���W�q�r{�;xS,蚸'r� V��C���)���?/�I��P`r	AKR,�� �J��@m��u:V��"�C����ҽ
��¾z^+RD"ii��g��1��=�㉿S�A�x�����,>�p���� ���>U������ػ���r�Z��oZ�q
U�$U��=��� 0���g����P�a�� �}y<'s��S�I�m���|u�.?��}�7�u;s��Jk�d��|�����M���
G(�+���g��6�7��������>o7�_�ݭM-�J�d�~ҙ(����}�@&�re��@�ۍ�T���@�z$�X�Jy��!sL��l��B�m^p�r�|��yJ��^�E�8%�4�d:*����A@?��@�+�m|z��E��R���w��@��⻇,U�F��a��C$"#9�������7lws�n�~����}���'L4�  � LZ#DK�,�$I�CsI`6��t8\��qaH� �����ý��|���rôX��+��%7��\�2��Ա]��{?h������B��\�(['psp�~�X���������qd�	�_"��p������֦�Z��k�r�\���?�g�{g��I?̩ $�&3
�I4^���,������
��HE�N�h/]�����/\y������c�ARb�?��d��k?�oH�l��֛᡿(p0]�{@͔S�@5��t?a���$�;Ɍ�׆6�W�ę����~�]{�3{%�j���;B��4R��+�A����͙M��7lwlwm���?��?���<\�^�aYlz������J?��S�dA�qCzy{%�~��P�� ���3�����=��z�x �X��B��^�C����D�Xܔ��L�&�NڙK��ڛ�"� ��\)�L^T�@ӌ(Z2(��d��b�狙%�6l�^���������}��Z_�7i9*iA�#�>p2E�X ˩�=�K%d&�`��"ϥ�] �+@��t\;X2ȸn��i�Qm>�v�=r]���C�>�ֈ��m�uC-h��ʘ�OO���S613k�Q)�H�7��Ch��"��>��e��(B�#7"~�����=�{ۖoݔ]E�`φ��H\�|��ѳt�ZW`�(�aS�i�&Uᰞ�U���m�]Ȍ�9��J�󟞿x����߿���*@�����k7_�P��[.�8�{:e���L��g�dBI-�a:�~!�n�v^��M&��+*�be�	ɛ ���5i�la/Y���9�p嚝�t�&��2������U����\g�|"�EG**�}6P�i��榽�ʋ���?o���[��>�\ �;=�"�����"�!:2�Q9�L1@���g,�I0A�Q�&2i�����l,</rZ'�QTC�'���Mo2G��:�����+ʯ��O�3_�u��d=ؘd�\O�hz��p��Wh�Hݫ�0�	�\���a;���}�޾c;��V�ٴ^�!9.�p8�O�=� �f��2�u�h���3@������|R�	p.A�<@j@^툘�k��_�Jfف�K1@P��P��GQ��~+�N����ʓOى�gd��+`*e%��ʽ����]�G��Nc/P�*P�1X}o�ܺaK7�[�Y���Mk�Z�ו�a��P7"UAA]4� ��.�[3�5�o+�%�%@˖������g�^{�w~ϻ_x��ݻ��������߸��O��;�� �ȞlQś�̗H���@�� �h
 ���!�Ky�ƥ�N�Җ-孟JX�Ҷ��X�<a�s6��M-���ؤe�����(á����ǆ�WSP�(��l��R��ำ���ܷ{��b��&b�H�V�"(8�f聅�E��}�\�Հ������u�̌����Z�1�LR�;�ێ?�\i�jG�66�5"!��z�(���xh3��
v��E{���5�?}�
����b�M/3>����4��X(�4�
��8>���Dr7-��/�h͝k�m���C�\y$Q�E�cp�vMV0/��Ȧ3��(�)�xz͡�N2st���p��z��s8�?�A���xXS��z8yO$,��%��Щʤ,[�\NY�X�.���3v��7�ً��2>%�S�A��RV�������ml#v��/Q�'%Z���ݿ���ܽe�A��[��߶n}�z�F��~�����Ǯ�j��}P쁽�2}.G�Ҹ##x�� ��s�M������]���c � �����n���\�@2C�^�ǁ�*���ǥ9����)@J���,�1h�����SY�b)˔������Hdl���$�Å3V��t�����7c��r���ぎ�f�t���E=ݼ�F�ۛv��f�ƞ�.���=��h�i��zӜ-*��(Y���k�{�ۃ~Qd2�
;�É-�@�!����ܸ����P��:��>����uA�OB�� ���*8&P�)ak1g�.^���E��NXy�*�l�4�w����o?�[J37�����e�{�e6�lЬ�����H����a���$gZq��B{ݞ)꽇�Z�G<`��8t9�Ʈ�`�y=��v�[�뀻�J����>o��	C�=4kS�#��4m"0�d���e�c6ⴝ<��O��|uT�$��(3���;h��5�S~o�8#E��֭լ���C{t��>�J6i�}�]7���i�f�zMZ\�dP�'����a'LN��&�%bԂ�8�F�9�JY�<3�'3g/|�;���W����������m�y��sݽ�H ��y�٣d�����r�dEܧ�+���qSc ]t����I.i�J��#EK��J�l����ج͟8c3'�Z�:a��؈�feL/�p詨��3�Nkh����Y�������(�0Rg���=��nYi�枭߿i���6:���1���p&p�*��|��R��2ڂF0@HK6u���.�N``�["  �P�%{X&�q���/f���
�.ƇO��s��@��ھ`�|N~�|�����*6{���N�Y�2*�r&����� ��F�!MTGR����$���������Ku��6���i���]	�v:>u.&���T��s<�{���!���3G�m�R��x��� ��X�'3����&��HV���ݟ����Hi�,ǰ���!bΩ�UF�lz�M�.Z�:�C%*̶X��B#[���fN�C��i'�ў-��8�v��5�^{dͽ)$��7�׬����[J��9��,�^cЕ�A�LZ��2�JU�: ��A0T�Y�X��ke~���\����{_|�2H�|>�+���͗?�i�+���K�gDz��@V0�2Hl��%���(w/�C����q�D&iIJ@�XU�^�h���62{�N_�b��Z2W��F׺=p��D&��4� �bƹ0��Z!�U�Wo��렛׮׭��e����7Wl$;��i;�w�`��5	�����9�|��C��	.UCd.��N��K���2Hm�p�V��Di��wȰ'���&��OF�p&B`�)�3H�֥q���,�aǇ`ݠ�ɵ�TF̊e�򖩌���i�W�,�.ZFj⮀�W�/K�(Fϊq�Cɯ,�C'`!��low�v֖m������Ys{�6V���%�Q��>�棒mB�x�tU�t�zDM��\��~4� ��D�Ka����]��cTL�T*��D.xKԊ��e�{?p�;��.��4?�V"D�L�
�q����败sK�˖��G�Z�糎m(��6*�k}A��E���0{��g�TA;�֫��h)m��-k�[wgÆ����P�n8nẆ[&��!&���4�vf�$ QMb]�H敋�(>m#�'~o������૏U�+����C7>�ɟ)Yc��ٳ̰/�6GE
�s�l, g��\@oj���)C�tg@#X�n�K���,���v+i�l��O���g.Z"[�� ����C?�4=�#.���ѐA���H�\P��۶d�f���e��V�x`��e��uZlV�E�y8 ��L��Sꀀ��������e������^����2�d�"P8�`;���WM�`�(
�"��	�$��H��,GQ<R��6i�){v_m������~���{�d�C@&e�u]s�̮k��}��)�s�L�C�f���NU�0�@�M(��M.�9�&�R���Q�B�$e��Fp�vz���)H��x�L'(�t��Sab�\#A�� %���=�(��P�17�C]02@f3���%с�&fD�GL�l6r���p����p]wЬP�J���iP��N�z��|&�c� �!A�����.�]� !(�
���f�]~�uQ*��y�5��D���m��0�D�����EDwa����n�1&�fvL�I�)9���f�n    IDAT|r� �F&�W�!E�@8W��11<!΋H�%@�Ca���!�ԃ�Be��n��Gdu��X���$���r<
��(�森ţz=/^�h�H���h*%1d;�( �D��ر�����������*�ċ������w~�K7$�v9�)NP?����<�'�*�
SFZ�͆���K�|_	c D6��@:sۺJ�b���|���Q�+IrB����F�Y���WX�������T 2���8�GmzL�I�׷-����au[Z=��Ey�'�nРz���*Km9�!��,#�'H }9�q#�E� W@���� Fb��I�x+8�� )aTl)�FS.��)@���:�R-G�*ф�	TD#g����O������0���4F�ھF������ųԷA��)�Sϲ��B*�f@^�`nN�Z���)�¸�������ըRmu��V����V�z�:9m�#�D Q4�C��-f�xpcOʑ�������K��������⸲��@$�G ��r�7q y٠�$�)� Q�@W:��Dk���4�G���)��?�Jc�|��hnj&�a�e �'
e�(�����UDC
)6Ͻ��"{�E�;�*G�v�B��A��Q!B��m�0@�r�N8�jL����� #v�hM
u,	�Ą=h]�Q������������~��ܿ� �x�����/�ϴ����"3p�$O3�M"�f5��O�;�'�����n_�#�Y�SPɁ��n��/�؞}T��#=] %�����p��1´��F=�S ���&��0��	�g��E�Y1p�4�z���x!<8�f�QZ�(�Z�W��~���U�|�\�(��5�p�Q��QP?�j8݋����ZWc�C�ɲ��t�h"Fn()�ʸ(�x��g�#E!�S���V�>ӊ���@�	����7���Q�22i��'%��^`P�<CO|ꏓ��P�k�e��ʤ���r=%x��FA��&; 4+V�v�FP"�^�Y����Q�fu���ł� �u�5j����t���.\B�Aj��\�`�-Z��ϣڢL�%`���P�;$�Cn�ʟ)E�9F�c���+�qC~q��GO�y"QX/��"���2i�2YR)J�G(S�d�LZ,�v�p��K>*a��L	.��\4�0qq�(��5�"�5��4kԩ��ݩ��(����D�_B6����h��A�	��F\@b��;I4bu�H~��#.�
QDƁ#3W
rSs�9�����X�u ��O��'����{�1���R]P}��`-��o���#];�)P�u�����wz1�&��:�)�')�/��CT��Cdf�7R�:u�H��5�(d�H-�
�HY9bdN��i>7!F��>�hΈ�V�
�2)��et�b~���)�X���ER=�\V�}�4S�H�(�:�m�1����'�IW@�F�'G{�d׵��17'"~^��D7�r�q�S�PO@y����~��,aB�v�d��2�x:�i]"_���>n��f�|=E��]D��8>5�m�P�����X�p����=G6����Bᩍ@d7������mҠ� ��2@��u�+ԫ�9��&n������ !R܎��rn�[�7{A�m��'�f4�|�]u�`e��s�Ȫ?��m��
��Q�udd&��ܲ���4� P4H�#MVɌ�)�/P�T&3[$3�%O1��5AF5�$G�bMa�����)���`�A4��)�( �����!��$��$r����d���C�pF�	�"qF���@�����T�xu�>�Tp�'/{ăĜ�'#7�-M�_���C�}�ϼtc����MO��_��#as�"�_#������W�q
��I�
³�k�}e��E!<2�4U��ƃ6v<EJ2G��4M�?L��y���J�B�|�����u`mZ)Ȕ���Q᚛\`ׅ)[W����s�&H�x�঒22�6�ǩv�(Y�}V�a.%����5W���#7� *�'��O��]/�(b'JS��KxY�2R�����k9�ceLB�E(�3; 1u������KzL�Q�8�5�(Q(Syj��q
�y&�}c�{��t�=��c�����A$�;"F�\1$×̼�\2 rз�?蒍�����>S{tBz��ݠ��j��py�!y|�ۦl�-�Y�Yrq�f���s�����I��J#�N$J���Jڏ��XW�ٷ��m��01~�0��0P�L#�.Q O:���%K���Tj|���������� ɯٖ Mޣ�)�"��.%����� ��&X��v�[5�/��i�G6�\�gPD-]�|�om9���|�X�'R�g����8^0���Kcǧ�����o�q��{��W��k����v�����׎�7�_3`�b�'��X�s����::���Y2"Ih��O�ذa:�f����&�����1�I��&ǃ��i5xkQ�f5���!2UBwO
70p2�%i��C��8@<񂺘jS"�Рv�*�n�~�4�~�T�aE��q�>ɑ�
ǺxT��<yPf��W<�+n|v�C$��x���n�Be]��2��	 �F�eH�8�ɣ�<�Y�\UMh�y�M�\��'܁�ly<F���G�)�%#Y�I�F��C��h�=��'fj H�D2��W6m���lq�q���ؚʈo��hRq��mPm�$U�OY�YR�+�.ed�h��!ld����N�_�	��)�#�!�0��ɝE
���ٜi�֗�]�/%IƗ�O�D�h�y�j�"C2�:� ��Lg(U�����2��y�U��Jp��<��B�;3iL���k��c>[�wd��E2ˑ& Qi>�r�ř��n��\'��ĵH�ߢ�϶E�㐦�Q�2�9)&#�n)�9E3�N��2�!܄�a'�|P�2�s�}]����;�xƯxT $�>G��?�X8�f��xD��:�;Q���E����M��p��&����<�mU� ̐�HQ����	*����2s��I��8bP0�l7���R�o 6�E��L�䃢��+w�Di ����i�(���.�*����P�v�bA�b��@!�`�¿Q�eaL)7j:�x��C�\VE������d{�) ��""�Z#�3�h�S�HR�co(��%_"���QBJ3�*�&@�����,���.��%-��v��&�;`�֥<f�������7�Wv�%�J�`�g�b���6 i*.�Z?� ����S�гH���;u��g����pAQ�a3U�#���l���B����۬]e�C�+�$��%�r��:�z���a\�(�Ȇt���u�L.O��iJO$JH3��	h��p	�y�Q\H�F�*Or�e6b����}#�"+[ԝ�͎�7�i)�ˍ�Ac����7P�l�:�5�`a4�1�*~O�!�S��'"S6M>�h�J�����9{���?�'~d�)�8ؕ �}�k7��V��U��~~�9yk�Ki�$|ϋa����Bw`���A�4���|Ϸ�T�ϙn^�I
�W2�܌Ɏ������09Oa<G��Bv�zGx��
 �����V�;-�SXm�� ���PV�b�0�X6�s{��|�kj����n�Ne�ʀbA�T�f����T�]��,���L��H4�;O�%"=u�Rz�k`�T���r�f#!� ܪI��%<X���.Y�3��ʳ�ATs4A�S!�����̥�
<���Og)��Li��9L$(��P�\�$3�${s�W�f�ɯ|S	�<RE&s�dM4v��]� HD%�M�oQ i�ie�Zz��.�;���ZEP,"V�L.Eu7V�Rz[]�6''l"�W	~���,R��I��3Ib�B���a[@F�m������B�<2u��q���`Oä\�@��=�������]�h:r� ��PÖ+�nv$��M�N�YZ�ŏ�3AZ�N�����ō�'��h������
9�6��E�h��" &����_h�J:[/�}F�5Go�H����ʏM~g�#��oW��9ʕ@��� �	�P��_>4Y[_�;e
�r����k��:�-$=�H�䚩��I�g��?�L��߾�߯����P�y��S��yz,ő:ֹ�$�'�Pnd��D�-A�+�>��QJ0.(	�R@�'8�uH!���;!:�S&0��
5�!\��8���7��r�VW��UI�*���dY��t��m�������P-|w0�`0U� �MNy9팈�g�O :r6V�)�v���k��S<�]�~�*����g2��m��Ds&�4)3�'��������4��%�D�D��Ђn�ybS�q':�XOhhn�����]�i�L��� 2�*b_%�8Tc\�A���D��uY�:�x���>���a� D7 ����v\4H�^ҦW�6��s�K#�m��� ���e8��@��-��DD���E���"%m����ġ׀t��d
9*D�w�<F��y�N]Hz�̳�cYP��(GE�D�t�"�t#������ܙF����RԜy�!��`��b��Sԩ.P��J� iv[�+�'H\@�� "dj8C[A�&L0�w@�R�*H?$Es������ا^r�{��y�ʹ�9�~$~����k�<U�����M�z���I������>pmv��O�l���R�j=�qzI�$�j5�ab��`Y�xv�b�7p��k�Yӓnq<y�Z˦L��"Eeez�&Y�bN��dE�6��l��M�u���v���)N���VS���o�ذ\'ce���e�D�7��6R��]�ڞ�f,�7�3i�qӮ��}?H������ˤ����M����v��8֨m�� p���a�A�;���V2�l�A�w\_1}-�N7E�-.�~��ۇLC1Si�
JdӤgSBLV��f$)ː�ȓn�(P�[1�}غ���)�A	�F�$0nH�RK��H�@&�e��h<{m������q��+dw��t7(t,�H� �/f��@�-e�4�?~� l�����1=@���聏�K#�5���Pap���@�PEL�����P������x����:N�ȋ���2D�Qv�M�(E][3(��R	 Y�%�����w��N*j~�����\7�[�3F��gwߥg9_��9I+�o��8�}�E��UjUNQ��ɰ*y���3�/�� �cXCLt�yS_�M����}�s�T+�LY���\�gs_��?���y��8�����z��n_lg����������<����k.�#��lj�Te��+�ɼ]vJ�B,��yd*�s:&����
('�Un�D��*�q"� ��C�J8�hr�u
��P���,: l���,��;R������GbF�n����%l5�s���f���f9��Ieݸ��z�� �[x���j~`�ILЩJ^"�z�����l�͎8u��9~�=OZ�,������3	��a�d�${���D�b�br>+��+8Y�cv�S?����-J��8JA�fK�R�=wW�Hq���7r��&�0�0$�<��nTx.�e"Y�qvH����wS���f,~_H���0�<7��]U5ۈ�=UӬ�sx�/_�t?_	CEa�MR]��]�3}
LE��@�M�<<5�s�D*�6Z�8��YY�<��X�)?p.dcK�DYS������0��|��Q�x��x��-�`�(4<1^-�Gxȵ�bADb%QD+/&i����j��<3�F8�<"�E��*���4�b��A��&��/B�@Qc�諊j.���n�V5M����N�Q��F- ������q;�BG�V.��<��W��[�A|�� Õ��b��/5����=�t��!��6 �IR�HM��耖�V�KIA��w!n�)\*�\Di+��Ѣb%h4\{R4��;���5���N/�0�cQ�����a�jq
��Ic�?��5�ЧS����=4��~�����3���_�;8��Fs�U���Ąj�[V��@�@�*~*Ⱦ�z[Bý��:��ó�<�8�ш�J."}� R�QN1Ty���	�VЮ-$�A*���z
�� s� a�����R��b6s�h=7��IN�D,H��g��m륶F�'
��岒���g��1�L���uJ�j��R�'����������k_�Z8��Onl������NM�pAa�TW7���	ҠnfH1���	����e��-o(l_OVŊt?y�)A��T.#H���bȚ&���fRh�ku(�z�z=r�Mr�>�N��e����z�&ә�r��"��n�L�kŭsM�y�g���ah,/n��x��9��yx��ǘ�����r� p�|4a��*�Ғ�/jeB�A�x GLo����4A�A���i4�:�NƷ/���K�<fE߈*Q:�&d�y� �ߩ������>���W�������կ�w����[��b6 e��i��P��Dl�7j^(?������df���=ґY��|��$G� ����q���4�y���MG�����E�8��'�T;�H��8>��#G~|��������/^]Yyw����� :��[+^_(G��X_̵�b9
�i*D�(�0���ሌ����	bH�![�lS�㇑���"k�"����S���&Pc����9f(�����X��T�]��l����g]��F��}z<��R[��Je�]�k���x��{'�@ĸ��i�L=t
��i�\74n"{��Miv%�4�f[�1�H�#��=6V)Рk�75jpH������}"�C$��$0F��3�̩��+.9��������ף�����j}�� pG`a���D35%���.$�.qy�(��b�H�C�*��#�H���\����4��c��rs	�m��х�+j#�a&����Zؖ-)�~����������z=��?}��}K�+��ب=�l�5��0YȌ����G��h�KD���l*�=�g\R���u�}ID�|O�N�h�l�LY�X�0��M(!jˣ���-��M�}�4&|c?�9JG�I��Y^����dr�]�x�3D��1�x<���^Nc�~���aRgU��֝��0w�"E��r�a{S�o�H�V��������=�Ȁ�} �����s�ږ��S������P>�Y���h�rd=Shs������U��_���z o���+���l�W�y^CD�%�1�f"b��G����P��(���M���=�t|�쮲���1L����O$�U���2&P@��ga���x"��B�����_\9�뻲�2��t���F��1>�&#_��-��RMt7�(~�&�����lb;_@Q��A2!C�����GyY�!Q��Ω�xx��e\�BRL������7U;��_�o��/>�i?sNG����q�X��N�9�n��N�=��L(�b���i��B��e@t��a��~B�W�bЙ�V.؀��nݸ��@4$�||�Am`~��F]h�Q������Y��T����u�6�f�ҙ��hi��s���}�����z��/��V�ٷzE�����GwP�a����l�sdI�؋c�Ѻ�&�>%���-iK�Z�%9�A)Ê��� �g|�TB��[�"�0��B��~$_�����~����~}�W�X�V��h4��H-Ͽ���Z�p���++\�1Ȩ����P����ZmHt��"$"���|���r~_��Y2:O�pM�8q�D5c~ߢ�uR�/���������w����?� r����^�ݎk���::̢(��9�����F�O"�9�:C�[n>�pg�'*d[p�2P�+'6��B�3ɦ�M��VHk��r$E"�a/�����Bs�;��3b�/��������u.7��],,\���r���%E�ę����h℻Ñ�2�[D*A�Ç��v� L!�6et�;�9	��g���$?��mPYC��<Ǎ��ϣ̱i��45QU�$�
œ�o��W�?��JjᵶZ��r�~M�Y���(_�^ʴ��I#.j�E j:O�D^�d��    IDAT�b�_�bBF$�Mf@���)�q�KB�W^D���^Y���f`d����)�]�1��1�H���(#�z�Եx<�6�|���5����q�ˍ�s��λ������]�P�7Q�1{ͤlt1!���H�"�sNqL���,C�ŉD��k��Z�ّm)T�M��U��	�9��Q�uGD�B�M�<[4fX6
 �j���6��&�94��㊲Ϳ�m�KK�PmT�cy�3-�%��Gb�-H¢�)��H!j��)�V�E[ym�曷���5>&@d��P�e<�.WH,V�@*�c�;Hz	��T*sk�X|���3w��%��5+a�쮯���h��o��h��G�[�p.n`v_hy"c�)�HtB�d�z�E��#�n�5i8߲��~5�߇��,m^4Xo�B�̺/���)9d��K$��*��z$J�����H������v�u<w�	�g���;ߔlބb���GQ���R0:��ʒ>. 2���:��9:7 � 9�HD-�ae�/�w����}��9�tБd�\��C�\��h�S��Mwld��޽�V�Zzn��3k�Z�9�w��D��#�x"I?�c cb�� �Q�:W�m*/��l?�X;	��SqA��������%�����:)/�vqAB�_#�%�^���~sd��¹��9������ʳ7�����I���^��;��&�CL�q4;�
[%���q^V)���[�_/�8�D���.�F��x���3K2!�{���a;�:����3ɫ/�>��G���Iy\d���َտ�v��b&7�xC��DWS(����n*[�D5����������F��QC�,'�/�e���i,F���> ��)�~Px@B��yj�e���np s<?�P��H�R��mF/��^7�<�����Wz��ի�h�Z �c}Fֳd"��ME⾘K�.+D�#:�������<�`x{�(�����D	�Y
��5��Av 2� ��B�D���A8��ذ*�`�A*:���o�Jc/�+���^���}����ԛ����?W<��&�9ys
	;�%���ɗ�#@n��E%������R�O��}-k�����#4Y#�mz�(a�M�B�R�:��UD6�H$�I�S�\<��ﾟu:����H,��z��\뵮����y��'FY���O���	4t�mN�qTZ�_� ���'�E�R`~T�6ߒB�T`�d�u�h� ����?D���rcr�1s�����#G�Ф�όq��43��u��u333� ׭�ޕz���n�Gp�1���@�#��F�{f��!�fMB��a��'�\K�
�5���o|��*b}e�zD'���VJ��1�)>��I�f@ɳ�ן��f���g�W͏��v.��]��Ƒz����^�b�� ��R��o)c�FJr���n|�K�ضz�&pI��m^?\?7Q�|��7t!9BgB=�T[��y��gA	(D��"j��N�R�t��>}����j�(<� ra�Y諝�����\ם����8}�sUMB?T]��� 0� 0m׍)�����bV�s���1l���1�w�\g�8�V(�Ȧ�1|R�\�BS6��P:� O�������iS���ITl�O������[7�<�L�Qt[Ӵ{���>�����W�ne|��zW{��%1j��
C�������p�6�	��@����<����m5�$��9J��t@��.ud��@��(��dl�f����|hc�8��d�l��k�F'�9����j�ot���������h|�Qm4����,<��q{Ð#jO4���mO�%���h��C�uŚlF�h�`:	M�t��2�r���_��g����N�T�����hL��rr��H���;W ����h4�0<�65EQ-����I��(���������)�#-����F��#���3���S׳ :x�x,��z���D:�t���,���:��1��2@�!h��`�����{;�n�oY���M_	u�u��b�f/�\����Z�Ca�����8��-Sӫ�X��G�#ux~~����_��l���Wv�ދ<�K g���F�J�-��rb�He% 	�!&B�bc��ez�L�d*'S<YO㳦nѧ���l�/#ر�,��/
n)~����]�j6���5*�疌�;j3��S�k.س�K���p��ju��ﾥ�i?��l��P0 ^q������5 F�a+�zQ�̄/�m���k� ~����:H�q�{3J���xrcF7K:�c�ȏ�<|�l�*d�"F�%��-�r�?&�����<w �����������e�W�k����A�T��}�Ɇ0��<����8Od)��Q2�a��Q;"�T
�d�>R(��v�/��=BX��~���@��!0)d��uu��4��=���ƣ���R��2T���u(�\jr,c������~x��������1\- ��������������:�&��iYUUu�^�#�4V�ٲ�8�.U�����r�j0�����l�� �WY��y��KL
:�\"��-p��ɔ�*�F,�9�ʽ�C�n�~�������������5����j��z�)�7�&�_���0��0tEEQ4M3L��E�,e�\����đ�m��7���T��z���S���66"�(E�W���/.8 ��pE�/ĐT�^�Ύ.v>��z)[���}���~/�� �Z5��7���;����S<��|6A��n�0;���Aʝ 3�#�LQ:[b�vU�1�2KC�`��+�|4�����7���=kkk��XX,o�����K�������rUok��'
�*iv��G��Y[�<��n?5�Hd$M4x���Ѻ�?���l�>��?KR����b�/�j�/��wm�*{�_03K��|�KA�0�0��~�q����yP_U�����8�a��n�g��G��;����y��l��=:�i�/��z�;�3�늪�����"���7U�kDU�uE	�m���Ov\��&�"I9$���¼FV��9�U�<3�׊��dd9����v��<����0EQq!��d����$�P��X�U_��n2�<���?�,'n�����h���|� ��ʜ����~ۭ���޻~��m�3�8�4�;����F�X�&V"=��x��Z}�
��b��09:��R�/I�|����y��!�� =��0�Atj����VI�?�'662����N/,��^�?�9����"F�l���O�7G��L��!��R��t6�&-a���Z:�R�	�c��i��tC�uײ5MU5�q5WqU/�}�0��o�N��T7�P�h�������ń�ei��*�f���*�g�n�4���o�Y?e���9�l���h�_2Jx)�:E4.(o�.���̓8��%�\vH&��a_St��|ϯ�>,!���B�\����p]/�͂n��	�a�u���x���g�R5}13oI%��^:?��
� �Á�P��[�}��o��U���TʠDL%SIр��KF,E��a�)�l:<���VFD8�����k���="M�G�Y��Xl����}���}�ݿ� F4��ѩ̓M^_��"qг�75=�'����K�s��h]W<�o;z����u�F��X'D�r���9�%�@��Xb�D:��N&�y�YH�dZ�
]���ѻ�V�ɤZ�Ř~P����>)�TJK躪)��6T/���X�Z���rg�T���o]��o}���Z>�)�2(���C��#��X�4-ŲS���B�đv')���h�x��/�+�sq�G�!F-s��;�{��w���Q��T�A�t;`�n6h$�uaztd��w��׏���Ȍr�9������q<�q������+z���¼N6w��i�q	c�"�����r9�<R~��D����>Z_�x^C�|��֛_|�-�|���r����F��Aq[w�&F�L�Rda�Z3)��5 ҈S&�����/>t��B��s�f>V~��0�/�s�UG������zZ�}L��	��vB3^����T
����X:t���?9����}.��ɓ'㋃��V�W��h��bSx��Fzܠ����mJJU�PhLLμz���'������b}� � ��[o~�mw������	���
FJ�3`��L�$3gdNJ @G 	k�\2OS�_���.e2����b��g��j���sy�w��u�^� )�ʢ&�?�"$�ݘ��MOM=p���l�k�����3@v_�����ju�9��eQحb����Ƃ.$�¤&�������􋞸���<^k����=ȝ2��[�}��w�����%6�1�,4f-V�e����f�l�w���%�j0q<�*�����/>r���0�ܾ�K�v��c��x�ѻ^

	��2�d��m�n8��*U��{jj����\q��ԭ��f�_����<V��bem�l4���R���rӄ+L���d3����K�ӓW=q�����?z�C��au*a����߼���o����P((�0y,�s�L�I�R�H@�(�4�\%�l��M�hbd��K�y�D.��ݾѶ�����������{�yN��tAzf�bD.�5���h���ANMOݵw���\8==,_l[�c�zv����]Y_}M��S��N4-#����)X�	&�hD�/"ä�����鹫.�w���};ȇ �{n��o�~��?8��`b��8��K%�:%�	1e�� ����B�QG y����d����ݾѶ���~������S�~ �f��W�΁Ç��фy���#u�3w�۳��#33w�vk�[Y9���J�����CD�2�f"7�7���@�]9���_�������k;ȝS������w�s�[7Z����؜©v&�D[v��
��C�AD���=��~kjdd���ۗy�ߟYXX�����O��=1��b@�L>8����BRΠə�[�߻�����Σ8�V*㋧N��֨�* R�dC�^���i%	�,&�(P� (�Riden~��?t��+�?��u�;�q�����}{�F��rf!��];�fӔ�f#���9�vr��� ��B��=3��G��h{���2̭���y�^Z��Ro��y�j�h�Dz�Q[��a�W� g��n�����<������o�/M/�X�~����wx �F.v������<��?bT�T*��ٻo���0|<h0.u���_>q�ԍk�ռ��T�T��X*ifr��qy.��?p��`�W(g�*狷�NL��Xv�bo_��`����f���fsCH�ٰ�uXdA4f�QvV�r5.#|||l�������=�����Z��WV�N-.�����)�,z]اÑP��Gr����7���(���s�{_���S���z�
`$���S�p����׫�"� 3ul ����@��6�ɡ|�s9��2����H&s�p��V���O7z�O���A�Hg���A�T��8D��Hxx����k���h�+�s{uo��0\ۭ�}mm~iaᣭ�Ə���R
�Ґ4���| HL� �,���3ӳ/|��a{A�bk�-��������Z-:�`У��2��4R(��Q�}>�![q��e�iʧ��/^���O�6�ÙV���N��_p�Q+�w{"�񄳣Th���/��_ta�FǾ<�g�����pm����y'?�l6����T�#O�HƖ�<�5v�jϑ���n�����}{�_p�ރ_��k;ȝR=z��O/�~g�Yg]HD9�@b�?�S�P`C��N@�n0@�S)7�L0�J�q,�^��m���s���g;�.�����r	`ġf�@��d���"T~J�������w��gl����>y�ӝN�0�q ��Ar��T�#�l��=�#�fL֔GG8�����ٳ�I�C�|������Z>}m��Kb���l���2�I�xSA�52(&��q �e��^:�����7
�ǔ���W�=����~�2��L��Ye>�3`!X��	ږ�3 �߇|�S���W��d*?���X���,.^�|��g�����5�)�X}�ґnC��x$�+�1����8�����߷��3{w=w�;�~��ɗW��o�	 �*(�D�r��}X���J}thDB�>F�X����ߚ*��?�(��7|�
4�po�V���8��~��4H��?�۬������]/�� ����'�K��Ld2��n��kkG���>�h�.@��XP|��������O!2�v�V@9�as�bq�޹��+/����ݾ�C�� �w�>�����뺃��C���I� A<I��Q�lN��Ͷx���0 �c�\6��C��ReW���� �z����\d9.d��x���󊎵L��F��Y�#�/��=Z�^^Y�L�Z��q���c��G�h� �����Y���h4���5�
�{&&�\q���-C���+���������7l�[�ݳz��:�W��B&J��K���g)�%S7��l����U#��j+T,�@�����ڮ� %@R���D���\{������*�+J���fk��y?~�}�ڡ���g���Ł�ǳȷa��0@��kA{���"~�����e����S{��Xx�?��8� wX�f�O_��_������C�nP���Є�$�Ѥ��2����+a&�c��w����(BNe��X��#�z�s�랇9v&+ۖh&Dl�2@F�� H�y�^��?X�^;��և˺�G����ꧻ��E H׶X�Գ0I�1@�:BhGRg G'�M�k���=�^d�;��N�O�:�'�^���#^Il��3�1�	�0%r� �dYNDx���(K����_4�� ���R�{������ۏ�$4��H%"�{�z��<h(�X,,f���d^?��5� ��w��_�h�?e[����w;,����Qҧ �Ll@��1N=F�l���+O�?"�����s�;��nw쁵���z�g��lt�j%bbcA��yd����8̰2��f�X|�%��0�3y�׻��h|���}�e�%.!�㩏� 	�V<�w
.��_��ޝ�d�8?d����-/_�lm|Ʊ�A�Ҡ�&߷����݄�l�yl��'F=�	&�HR>��mlj�WO��z�!@� ��^obqe��^����?wO]�^6ua�P��p*��K��'��Z1�}���?�� ��>�4ױ��
�W<���5]8�z��� i��b����;J%�t�G� ��F�v��v�\�U�T�I��,����	%OP{�q�� Y*�n��������;�v@��_Y[�T��}�a�A��Ȳ���@�mIC�Tx�銡̲�M�-e�W��7�vU泗x��{�z�v�{�'�� A�Y�K��|�5Xg�jB�_.��T��xϸ�<b��F�sq��jk���N�P��"CSHgGN���mtU1a��6�`���,���63����cc�~l�;��v��:y���N��!g��qBD� H�6Þ� 1�}���f���"���ө�9���d۳�x��R�V���{�$��Z"W!V!�\�#�T�q��z{vz��Z����!���=�n�w���Ϯ��]l*d8�2�d�T�]� ����KQ�X��ٱ���^z4^��9r��F{� ��,�x�}�I���'}��8^�Q�S��\��)��M��_.��P���5^n���V����Y��� ���C1R�c��#M�? �- �h왜y����ǆ�3�x�u��|veu�RU	�T�1@"2G[Z�)Ĉ=�׾��1*_�(M�ڡ�ٕs	F���5ȇ ȥ��O5��g�ƈT^)Bee1!s�P�ߎ#�@@��g���>��cW�$���5^�t~t�R���:ӶT�h!$�	��f�M����H�5� �{�f_9?Z������Z�O�x����KѤ�gӤ�0� )� Ŗ�6G�����r�P(|i�4q� �z�;-��?�h��*O�lHNV"��a� ���̦ҔJ%������Џ��E>�l�D�V��㹓����'ll�57  IDATG1�5GP~T�Bp�!!�4E#]�����������E�����j�੕㟫�W/@��B�A<1�~�,]x�݂����@\��A�b�oƧF�><:��ۗuA>D���xS���qR�bo�o�2;¦ !f�L&�L���S�]O�={��5�?[�6>��ޘ�QC��qqX,��5��KJ5�llJue/;89���~��~����_������f� )>
�f��� ���و�]{�b?��R������*TC��ᄁ(�xz��n�,e�g ��i )(p�]X���I�A�R������w=U��%�����Z��n�u��N�'\��W�7���"�B�t!d�A[]ٿg�KL��� �\�;VV�m�g �_��cG��T�h�MU�v)�G�޳����ҢVEծڵ�1�R+FK�*�w�7����>��y���s��~�S׉�ҼJ&(YVY��C�N[B�3�`vM�PP�ϼ�\��ߠ������%x����r�r�]d���=��ҭɣ$>S��q3�<p���veh���T�����6�>?a�ԈVw�t�~@�پ�ʳ}��_���fK��!]�uW/�������[���/���"!~�XT��n�brН��J�I�v����Ɯ��>v�2�DT>��N!� �r�v�x���b��J��6�hˡ�[�KJ�ut�M��lD���+��I��P�z�}�j�w� ��Z���*w���2���a`�l*��'����J�kf <���P�����G���6���,��{NN�Ƽ���)?�6��I�id�c^`t��]M���]���1\����s/
e�ڰq*��Jɭ�B��f|�fgTIL�hѮX=��������#��ȧ���Ow0Z+mE��9�������	�g�E��5$�D1�i����4Ⱦ�:���3r]>S>��r{���+�{��U;G�f��<4��y�y�fDAW���dH	8T����t����䣠Pū�x5�o�ٻݟ��(�6ˌQ�p#2>\�'D��Y	�a���_�88O>L����lu��LC�3���Y&A�q�Y/���X��҂5�Ah��+���ES�(g µ����8�D d�[d�z�Pۯ�W>&ʹr!��Ř�ϟ�+<����������{Ka�y5���ZJ��_��/ܹi��()����G���>7.o+*���Q������H=��1�H��%��w��FK^���b��ᩫ�k=�z�Vf�B��=����Am_�6US�
�]Hh?N�����d�v�=�������Py�z�`��x���d|�>X���`(0Idq���� ����tD�-okv�î���D��a�J 9�z�/V���u�-���Y���ġ���#Y���<�Z�_bR�kj��J`���~_Ĝ	..j/�Y�8ъ���!KL�����:���e��hp�Ho��Z$4ZR�����c,BĈe r��G<�J�>��?��X��9}81��^���$d��N*����̟d�@��Y��Ɣ�U����wz%~4����ө��SU@��B>@ O��NfDd�7i�hH�0��S��P�@^iA��9��/���	V�ζ�SlT��^å��>�A���{47��~1��/�)2���0/�_,��6K5��s����� &�<hT	AN���՗.��Q�3��YT�m��BYzY���?T�]iT� $��7L��#��Yi���������cݵ�b��0~ˋ��-�oUƚ�r��e�5�ͼ��}<љ������B�x�z��g�U��3C�x�aa���Ņux��[�J-��U�'�E���6×�T�޶�)�
�|���`���t:�iLZ6�l�9_oM�����F�L��h���8Q��h���V��������.�QxU�y��:\Dz�������3S�_��b�< 1n�l�GY!�q�87��������	����i�Mk��4������ K}������U�a�P~�Ç����5;s ˶ ���>�N�_+ӷ8zkjV�M���3���E�&Ϧ�GZ3�������Ú��7���ۆT�^Y��~��Ý4��B3U&�/P��݋)f���L,�2�ny�t�\��%��9~ni=��h���7G8����;&q�v-n��.���26��n��=�n0A���"V�XiR������<Sp���#�UN�6%�Z�M�@���{��s$�}{4�ǘ��K���W��ͦz��zV�s��� �e�޳������I��I�_I++�lf��>K���!���w�Uv�]�����8:,yt�3��=�@����o�n%����Eܜ�y�E:���Umy�S��@t�3���jJ��}������l7�y��&��7��<���G��?C}Jͣ�^!r׉v����$e�E�e���r�hG�q�?��*>�l��W����g��Hw��<r7��c�˓��(�K2}a�DG��H�2V�jƞJ-׬H��N��=�	P���M��Y<;-%��4:�v���^�/7p@�
�eꃹ���KMbS�\��T^���8�f�y�M� ӝ=A#�N��R�o�C�Q���ӜW�̉-����?��ͣ3�f<q�@�];e�v+��B��e�����>5���a�$
@�˭�u������G�;W�h��d�o䢔���Vx"��͗���kh&��Î9���x`�d.�9������A��r>�/2�_�e�υb����Z�o��-�{4ES��^t�~͖��XoM����
���<�=�WNm�]"�����[��5�w�K ic�C��U���A_�ۄ�4�dV���g<n�D]���f���Y�)�N��:r��:���8��G�/4kt�-��s�G�|<��C=I����Ms��PZ�Sᄪ���Z7��)�:R��U�N�wo�jzd:Y�2	A�-υc�e�)w64���T�w��׉����~�yR,���!�M���6Q^�R�d5�Ƃ;P�ߎ�a3T�%CV;qMЕ�WXȁ{�JH�jz}jYN�{2���Ͽ5�۲����5ᮢ���V��œ�� @"Etf�e#����	�r1|"#�Q��p[C^!�a�JĒB��E�Q��9q�u��i�ɔѫO�ku��w؆�h�����������?m���E�n~٤�R�n�%Ng7 �d��>�_9��*%{g�
{�Ƥ��?i�Nm�jڰ�Ӥ�~ɣ%2�c*mT������m	��U\��7�qF�A�N��<�α��j�����~�����= ��T�����A����9�7�
��q��!ΫH^F����L�FA��8 ���M{��](xy�%�S�У��&���O�n8��g���4��(����8XQ���bE-p��V���j�J$�h�1#�����W�2.R��G�t���m�$+���qu�/ڂ�S��5h�^�u��r��N��)���Pq��lݩx.��%|&:.(�"i��N�b�+4�ӱ|84dk��p5��D����|"�6��m��J��w�M~�v8��z��P�{�9��W�8t�O_^�@駛��|����Ӊ�ǐ�t�����?�?���(7���!����i�ݕ���P�9 .��	�w5{]hQ[� �_�m�����`�aئx9˾�:�>��n�����m��mj�z�����EG��3Q��ߛ]?ȯxtZ+��v�sf)Aϲ�U?\�oy	&h�Ѽ�J@`����}�Q���f �7���O O2 ��O�\�%s�g�
�˙��ӲF�[C��6�̱Y�	4�8a�2�'=�|3_�p�F��W�N�@�#~���-�*+��z�	��j���]�m�$����^>��7��)��$VE��y��� �@v��b�OjJ����X���ϝ3��Q�?�O�����i��		 ����H�
ִ>T�pض�l�g�D֋١~��W�pZ�f	�ji�u��Rȇ���� ��g"�|R����[�2�WDdT���S&RYl�
!���^[R1��}<�8m�׃�F3�.Ǿp�_*����O_�m[�kͧ-�!Q�f���YXd�5�/��s�5G��Nt�����į���j���c���j�C	���v7�=���7QY�Ġ@�ӓI�< �����sd���?�b/��,����;|�}� ��Q7����A�BH���ݽ��i����a�>���Z��:����j�q�$\��aJh��gEAT�nŒ|1�r�f��\�������:ۭL�f�s��V������*M��_�p���� �C_߰�G����r/��"�SX�q�tZuMWP���SW�q�	V�Ҷ��SF�/,{R�=DZ�
0�׿�-(���=�;?߄M�`�'(_�t뤁̦W�=S�|�9�j�R̜����oؙ�i
sf����f6�XBdw�Z���/�Q��V	��)�CؐE���}��.C�&��T�k�=
� ��J�թ8�	ÖI�b��[�]O#���U�P�	s ��4��R�A����X>'�m�
~{>��k�Q��
��C�li�fm���pN�F#�\�Yk�������]���iK�������Eh�d!��u�_�D�-�1�&�OŤ��
߀�� �&��[���Az�>��Kl���x̯�T{��� ��K�Z�i#@���̎��mǛ���2�f�`W�!�8�����uzg��]^Ȓ�狝浨\��3�\ޚ
q�ؔ�	����Ѧ^,�W@�N�Ѐ�R#ߥ�x�u���o�/.������sCX�^�����d��9�)�*���M�NN�ݸ�d��Ξ��K	�]�͘�J�y��Lu�E@�O���g��|w�'VȽă���$���*��s��7�5s.>؊Vl�R���il#%Kq� �>$��9�!K|�n#8���H�A�A�r��e�E�����_9�F�{_��y��������h���FbDi���5d*ֵ]�RV:��v����R=Al��P|$0��{��<V]��m����<�*�ԛ�\$oB֝�Q=db�BI�ONb��;;�j�8{�	䈒�;��ZY��OD�;fQ��t�=mA�.||��FF�}���ē��C�Cl@Ǒ���3^M,�QDcO��_&��/���:� #7�o��6����[�*�.\E���K�*��2������s��by�ߘ�60u���w�����
�1�s��O[�L<��l��^M;r7:F����͊��q��{	�&����ҷ��+|��Q9��া{>A�V=%���N1�r�:8褳=�I��,d�ZN�	������s��n�[�g�ݟ~��l&��I����]��5�Z`zh�VQ��^i�p[�tZ��&|�'��\w�cڅ�B� �~�w��)�ͣ|��_��V��C�ø�ԣ��
�֣��wOVQ|�E��(1 �p����Z��@��S�]�=��?��-L͞g���(���t�xz飼����;�gH�ˊ_�K��RM��G$�������lL��&�R�yGd´���^��tMMK^����;6�q�Bqd��@3m�3��a2ui�����2W�S���%jv 5�}K�U��i���������42�ƅ�d�B���W�De*:��u�r���^2��g{u����m�ҷ>�ǰAħm�][�Q(#'C��b����XƏ'h��K�1�H���ە�wh���^���w�^f�A)l�E��%�'C*ƪ�f ˄�R��`ќ"�6�����[��={NO_饟�-Hf�W���5I��[d���+�+~�7�7_ÿ�)?W�b�B��Q��,OmN*��U�?Д�����L�(���Q�$��3eݷ��п�����{�����ŭ/����u��b��,eO(�mנ����#�aǮ���>��
��7+�=q�����.�:���.B#�YSͯ��E�U�|Bh"5Yu���K�)�Y�<���T��^ �5?{�-�`�N݌NBǐ	�cdi��>j�EkO��ɨP���h'��ٹY��C)�J~�_=�v)~�]}�9��dc����y=`��=�Zt�!�]Qm��7.C��Sa5�>o�y���R?�����+d�}D���N��g�{{��1a,��������U�$YV�Ô�E&Q�vN�+t���_���݋.v�o+�Csy��8�A�8�!����F��R�e�n՜m�6�(�n4�T喕|Z�k�s0��J��t�!ne�����[z�w�Q�hL��>��LF����|����H;	k���ϭO��"#���:TQ�i���v��ǲ��e�_�Wr�O?�����0�6zc[�n��A ׳\-tq+� &իɡ��ã칔)&}OLl쪋����G[��=��E���z�os�+�� ��V������.���sN'G��S<%^0�@!]Wò\r]u7�@oB��2��L�f�I���� $S�<^�_A����g@RⒻů����:\�n�4U �@/�~@��(� �Ш�|׭�%����_A���ïX.&
�?O55j�b�PK   �-XS��
�M 2T /   images/a053b5f3-ee57-4c4b-b9e3-486563af4e78.png�{cse�卍N�۶��ƶm���6;NǶ:vұm�8��L�U���éS�k9[k���D*�K"���  $i)1e  ����eby;���EYRP;�w
 �ńU=�/�-���(<�u�d_h
*E��<�
��c�V���c��DYH�Y��Z��&&���/�/��	�V\��{R		R�HٗRMP��7[���"/uҍNwK�!x���"����+��&|A.w9ר����H���Մ�o�?Hs���l�p�����ca�����ۡӁ� �?f��8������t
!.h.s<È��.�d/E�j�);k��§$!���L�c��WC��
 a����EJ�7y�a�������P�n1�Y�Η�Z��!��1q�~/=P���l�z�t0�e0�%E�ZH�hF�O�,TB� ��7;���[�R���Bv=#�f�U��o&fS�F^ DRh��O�3���\,?�uID6�|h��{hW8J���Υ�O�r���u<N��m'8��	B����F���1?L)pO"yAW��U��C�5���8�@��!�`A�9aJ,����Pٜ-qn�D���N���dN	H	,
E�ϥ�f]Bl��S�������P�K�����)
c`��&W��5�ː�8$�qU��cu�lx0��s�Z'L�wQ|;�]KK�[�N��x��C{����o��6+�2�H���q��j�>��%�{��갶D[��R:;���FZ�-��5��*�X$\L��䉋�j�&�/ ��=kOU��(m�Z��e�"��o��|����bΏ�&x�I~�����e���NHS��0�9H4M5teH�`!af�6މ�O�8��A��:��L[��er�e�����u�_�m��?QE�	F�G������<K7�MM�Y$���+Y����j���9�ZjZ#h��5O�@	���D�G�Q郰�SGʤ��H�`�*^x����(j�9{V�3�AF#��h����k�i�toG��(�E��
!����aw���E?�tM�����<��*J ��K*I��;\�^'�w�*��q�EGE��R,����~cȜ�g��������]�!B}���Ѽ�ue�r��[�Z���4���;5fg/��]�r���c(4��	>)
���F���)����.�
�sm�v:�2��eI�*����dVe��h8����#K]A�!��?6i|� ۭ�o��u2�k��c(vd�7+m��o*�x�B�P��2P|��̬�Ґ�a)'��F$��tN�Ҧr����Q�;$�xȶ�<��#M�E��_9���������L>�����a��1Y+7#s��z����Q5��M�K�Ss�֪��e,����TK����L��&��p)alZ4�yք��{��,��
bˠ^�}�gLj�1��8����͊⎣.#���:��=?W�������=���p��-�9@}�WO���C�܌��	T������t�f��M�jι�y�CN{(��4�ԔF�:�B��;���v-�L���>����r�5�Y,XM����g��YoNڋs���)L�Q�c�_+�����]�2V�U$���<%q�;�H�A�j:3���Z��4��u�CҤ����S��L"W����Sp��߳���|�Eɬ~�%����+�N˼��{���/H�;H�Q,K��e�.n��#N��>��,��8⍶�2�\AϹL��p
�tN{bQ�ӱQ�	��)nGd����s��b�u�v�' �C����NsEn���%:���D��,���j�O�#��=�����ؓ����V�O�o�$�UJ�7��D[>�I%v����9Nz����	9�.q.8Y3��	87�J7�B�����o�!�A�>1ץ�_[��m";������[����m �ۨ��Ӥf�h�Ng�H����V�* G�q )����s�$�#��H@j��	�e-��% ���s^�N��V\�;	7��'���6˅-�+p00Å��nHѣ@e�~�X�H��-+9�-��h�L�uXY��>6��p	��TB"�ы��H����֧", ���0cNY7�2���H�P-t�q��#Z�D��p֗��'(��z�����U�1�#���
/zW�4/��zS�I��<����n�_�9ɾ�����4K��>v�Ne�X=*��R;X�ϔ�S�G�"QZ�T7P�D��h�2�Şe]1g$�1!e�W�z����AAWl��#gv�������CoF�ٕ�&T+`���~DVd�����WF�(��gw_;��s��DV�й'	}a��!�X!>�,�QK
[����ռ����<�♭L����R�?A�3P��('�k-9�#ޠ������O��:ĺ����(#ʰR����ا����PL�.�#��y������N����Pؾh�9ce�=�č�YZ���(Ħ�b�GM�WR�DZMQ,��Bq	i�G/���I-�1����V����"Q%�
,m����HF-+)˚�����6�LQ��1�g�������w�¯���Gx��qe�I�h}��;�4�T����ϣ�Y�I��/L����,��.��-ؽ��!�($44ׅ�Ũ��I�]n����������$q�,�Lbږ�������`�ߔ�1��$�<z����G�������׬��­Եu���8a���2Ӯ�MZ
ܰ�]��PimJ���他�.#TƎ���]M�:�j�T�n> ����BF*�$RM�"�������As���MD@�>o��3����ٴ��2�=�s}�`묜~��q�6"o?~l���)��?��](��>0Q���s��Hl���-�����ǖ=�.�=I��I��;RJT)N��5��):�rb�kLTI�F4�W�� �M��=j�\��g�X�&��)f8�ԡ��	9>�н�c�dj����t����`��|��������f�j�� 	/N�zB�ĳ�m{���US�V�[yȣ�lМ8�j7q����;���I#%Wj�1k�7���N�]��i� �J�d
�^&𘣏ZMF�,���E�F�'��N�Qx!͐k=�z��Ę�+9N�\��֕�L�wMa�RT?��Ԥ��r����	?�r��XK�,����paf�xL��$m�׭�NR�g�����6��~X�ĝ�� +�]='�|�-'�,*wiU32	���A:�T<�v~X��2�9*N fj6J�����ד���w��wG&��?��m��`���[����"�m$���6xx��/��\����q��W� z��G�?�vx��a�en���s;�Y�YXP�6��y�
աE<x����e�����\+�ڂ���Ԭ��ޗNi���Nh`w�)}��2�h���['n��S��G=��"^R�I� Ԣ��;��*�=JX��%4�S4�׮5�+���%&�����Bo �B8�f���c쉔�*�N2ng�UM?�z���Jw�nu4#�f�s�ڍq���үTi��v���p���	�p�Q!��������s��s����/vA]��>�lx(���Z��/MV�S�e7O&s�*-��<�H�`^�˽��uz���[�`�$�.L�0/ξR�YVPZ��s?_�
O�D���x�ړ;{j�!?�_*�%f #b�;�t�Gt�pS;�@�5m�aq���iϔ�pH����$�t_7��p�����Pٺxl��c��|f�O��Ə-�lO�Z����C=����v��1z�}���>�����9(̋Y� �=��.�O�����K��KϕFV:�Wi�áY�����Mw��-$]!���V���h�b;iizxڌv��ܤ�d��Mc��4������͙����F��J�"�Ĝ^��A��C�B��(�[YV�al�j�t!u�;eO�SD�B�2���t��µe�C]�f7��v��:�f�ˌF��W������
Y�ӭf�k����w�y�ʥ.���(C'�����\��qs���ؘ�+{�LdJFk�.��8����A��oU�2����v��U�IK��)��l.�0�ӍM&v�OV�z���l�BV�{����ݔF�y�rq	;@(d	�Q�.��(�m���dq`�X~���$*Pچq���6X�Ӝ��,x�<ɝ���LH��X�i�1�SɁ�'�h��t�����W���K?	�뭩-,�Q́L��M����ؤ�c/Q���r�RI��ɉ	b����w�N�,��̗��G���� @]�Q5�a�~�·Mg���%���{�֣a���u(�A��.�k���p���&���o��qͲ�\KN~7gY�'Ϥ���*F�9R��Pq�A�X���P����{d�J�\qı��:���e�]���d�WQ"@K��O�̳ݤp����߶G�-���Aә���o�+Տ`�7A����}=~gj^��!ev���Şʹ�����6wԅ<r��b�x(�m;�L��*���咁ݣ�F�]S �48��S�Y�DW����T_b\���Xңz�鉇�X ο����yB{�����zY�>��5Ͻ%���ˎ_������h��'�h��Kg�Y�;��,a����TĐѦ���7+�U�
��l�ҫxwwuxF�g6�W|Z�V���l��T��,!�g��}��$�nڸ��{�xjȟ�y�C�[��E( �p5�����#��n�PXP;�,\v\VBGML�B��ё�FT1����=��:-�@:���'?�,ۺ�G�^/7�Z_���n�3��q�j�?-n�<��ӽ���+@�L*f�|�e4��[�L/,��Xcc.��v�%�Yi��*�zR��au�MJ����w�g3�gy��]Y��q��>\����{𠷓��W$���~��9�x:k��Z�qD�rHR��}��`�Ȃ�pC�!`�D$t�y؜��!��;,���ˑ-Y*_I<���z�гY֭w�p�e���aם��a���+(��k5���v=z�:*u�	�E�(2З
��ǲ�-�ŉJ__WL�^<��T�� fe�<�+��[0'�"�u;B�����A�޲�7�7Q�j��� lۺ��"i�r�2c��]��if�ff��ԛb;�@�_"�ׁ���[��0��P|��X�y(¨X`������
��}1�9���!��ٵ��<5�<��.���^���vr#������N�jJ�݁�S�Bss���OO���_�ŦTG8�޸h�uԞ�բT��Ђ�ON�9���##�Oؕ�8#x5��e�L�\�X���22��WXI�S�jե�ޯ�Vs����'�&�c�����O����w1�o,��H��u�k�Jͱ�������^!"\��\�H?��!Bo�L���v���}�`lu��
�n^�%�S���h��}Iny�],��HN�d�|:�3��6(�v/.�W����cJuF�KSFN\ب���U�d[�*���V������0_<�TLA�����=�X��N[��]��`���Z�n
Xn8=l]�`�{�8=U8L>�Pd`��=5T@e�"HL��?��I0>ųc�k�\|���.���
^�J���,%�c}�����»l@tnw�a��%pW�-���s�+h ��E.��ao��>?j��p��ӌ��Ϋ0PΑ<�D�,�X�����ēEUPE�)��	��p��,"�T��c�O�f�����p"�u�U�7�^�dx���s�_1vI��0諡~6L���3�����QG�YpD�,܁F��Dl���~�4�\�^�_B�
����c���?��۳�d{���g�����0�Ņ=�ܲ���t4|�|ѫ����^$K#/�^��,#�e�
�9ǚ
S�r�x�K�ܾ�f;-�޾W�x�O�K����9�j7�6���H��Bf�#�w���.�ػ!����$K�a�1���x��td%���N�~>�E'H�%�܃���f�"���i7>)4��C����j���^�yӷn0���6�؇	��3�}����� 7�{^�T�$��)s���H𻹖"�"9a{P���ȒGC�k.��uͦ��Q0�=�>�p��:����=���o�tt\��}TI�}S�9&�_Âa�y������/��bK���0쓜:+��j�[�?�E|߂����eJ#��U�a=ЗEc]��b�`�lՆI�M9��j�on��?�m���OJ+�$m��	�^�}-�����#�NC�S ^[�F]!�P�<���M�g�|'Ͳ@	����\�w�i���80�������ˬ`�g/������� ��>܀���ѭ�l<<�I̽~���rB,�7���`��"*'�MB'`S^� ���Q�t^"t�C��$E��gϵ5_�����R�j�6��T�g��ct_<���(�`��o���Y-���~�ˤ
g�#���X��
��eIG��44*D�!��s�������4����42�f��ll�l>2��s���Z�H`h��
dU�K��v\IM���������7M�?��+!�"�`�N����C�H{ai�r'����O���ͽ������7���1�O���Y*(K
��O�t�vX<EΌEV��Z��U'��P��I`D�L*�֬�������5c/�
��U�w5x0�	|�][V۝W�zu��E�E���mv6R���\����S�~y#0��heN�k����W >�y�lI?�{�Q������G�'�d�%�#ә�,K���~y�e\�kG������:.��B��$��FZh�x�L�]����ʰ`�!�R�U�W�K�"�Y��-`Tep�� �Y�����T��F�|��)8|�-K���Z^Ӂs��Y�{v�=�ߌr���9����]I 5���'���l��k�ΘN�Z�,�1:�IjjP�g�$\Z}��{�go�6�� Z�/v�����/�9IW�B��9�6y}����N��K�}K�J�h�V!w�Ku��h,���WO�o�x����Q�pԸz��Y(�8ެ'*���N�G�����p�؈������,27���D�]�¥x��>�H�+�]��s;"d;� ��G������ZA	y�Y�$���eO�N��f�1d#����o�JFE����	�׶e���'o��.��
��)I{��m�bI�7aE&�̤o;�|��Dpm���zT�%3�nϺ��h����
O[n�[��+��:2�]P1 �c� ��?�.(�N��K��.�fr�?S�9'�d����� ��U�I#���CU~�A���W�~��hؽ��;$��\���_}��ۤ�bj�o��B�+�hg.�W6*�f����ղ�cu���j�SH�����W��0�ʈ,I}R�T\�d����V�)/��i��g>�U���[{H�	QߜW_�y�.��~���[���!C|r2��-��N;�{`� u� "Q�{�gӁҡ�b��������K�p6Ǉܺ��^�˹������J��mC����1Z�����?�`��0�����Ǎ�%����&�$H&(9x��E�`ނ
�
�Ԍ�A3A��u����4_ߜ���{�fl����[Zl��}��_ɔ���r=-�8��X��E�,��<8yJռ߃?A�P,��6I��qA�{���F��i{��=�b�j�����z���D�K�����dΤW��`��{2M�N-^������}���]����,E8,�}��c�{���u���ya$��Ix	k��(�o�����k-��ؿgЉ�r�1v]ƀ��e�E��δA��sԮD�),*�%�Z�P�l�]�h��{�DJ����^%��'�o+�V�����M�/�zv�DKڛA;�{jʜ�!��@��M�w?&K�\��D���R���7f9�2}�|t��a�Qr�6G(���l�����G��ai�D��̠Xˑ���)��_�r� W-�9�I�D��#u��1�Ui�����M�r�͌����u���^*�+�\w5|�\�3�g��w�����ҽ�J�^�2�j��A#J�j(��VA7�f�E(��W�!��9+��k��]��+z��j�8��:L�+��"x����Ρ��Kw�Ju�|���\�W��o��N�(v(�w�q zǩ�����D$��O���aܛ>9
����r������wg�tV��D�Bn��4�K�a��IH��TP�I-��^��K19oN��2ɁE	tRd���@>1�5���z?�Dヶ�t �%!���@�?x������M}oaH�Ŝ��dK֤�j�N�5��E�m�R.,�R̄�P���s��x�Z����6\�k�y�+	m�]ya�!����\^���e2h�%��4L���E+K�~�V��'YC2�a��c��R���Ki��� ?[����Q��`р�٭�~Z�^ϫ�a�V̉���,�wIOe�����l�(\��1P�w�c�}��D������I��B��(n���ֿ�����%q�xt3�����̙�>��2��fˬ�g(ύE#+zv�D��V밅.-�-\:��+]3�L�.�鼾p�լg����o�$�m/^�~�wB��Q���������R��ū #�);�)�s�9�}�\���QKf�x��=���a���q"�cZ��A��m�}|���\�O����D��M���UJ�P�A���)�텧%��i*O���C�0��]�ZZyYͥ�mo�|�	;o��<�+`���ʦ}���
F�'�������+T��Fk�C	)�(�+`D%0W�87��GOP���D����nߒ��LF��
DgD�M�}�s�@�m�����JE%�j		q���v��7�����3�����l�Vԋ8͔�3O�kaǸ?�(P�BK�)u��	s4�y���G�A�ׯ�ӫ��ϖ{�1kn_O�6�ZS8�!IGB����ϧ���v�^�n�G�ve��
nSSx�H�E�����ڬ�L&e�����i���H�6,o�f���Bޕj��k�v�ϗ��\WI	��On�d��=U���O��&���=�2;��.U�$61�XE4 1�B��B��(E1�HĢ9�P�����Lqk��FfW�A�Q�CY&�̧�hC%�s��� a�}�8��LG�ִ���_|�;�-+=�䊺�����T�ku�HB���8���?�o�OU�_��g,T�,ʺQդ�<���Â�iV�W��򒑱v)v�ń�X�(��|�Ñ�z���"�ά���!��%r�\T,����x}�.:������Q"�V��mR�T�e��4f�y(�(F@���*�(��T&�$�_��	�W�[�AWm��j�(c�D��C+�El�#��*��V��I��.%�CĊ���̴0�v�*��c�b �N|��zK߄�ߊS����^�-=��v�v���f745�CU�0�*�*�Ěƫ���ҕVP�c�rMb0��{��}+�|�n��["ut.��du��=���A�l��Ku�o�x:��~y
��.���[�P~�T�`��P�ڬ}.'9��LxX�Y4�"�Y*E���ٜ�ݏ��3��
�2��G�IDa����5��ڣ����`D��-OP�W��Rb
>��\x�KzǐB���?P�*kg+�a�@��l�s����]�s���N]r�J��Ee���y�����IIUO��
iS:�M�%ǥ�!��4%�7�d\�r�����^��� ���lV *lY��0�\�L&x�^��./A�1������L�����) �[��K�ϧR��H��b��w�Q@������~侫�W�����C�T�_�۝*>��F]*~�౽��q��/��X�+P-��y1�z�Y��C ���	�u�e9}$�9��,a$A��9�ty
�^�t�~����b�r}e��
�6됚�Mx�Bȅ��};�j#�U˪�]����K�B�JTN)�HK
�:'0�<�XX$*�v�����%z �[�i~8�Bp��~�Be�fSw��h^\��S��fG�d&���HSICf��Mc{�#�Ƕ�,����J-K��|�q�Z��"���K�ՃG��	��R4\d�(N��Z���b{�Y�aգy�!Ǐδ���a���F��� �w�^?�u������l9ڢ�cT.�l����	J�u^��n����s>h������Zl��n�Keҋ&��]��w�Z=��,X�m�� ��C��K����B�M�	���
Q0��S2#�dae%���������{��O��Zy���Ck�����>��Y>�͟FLK�d�as���e�r@�i�����5�eB�ɹ�c"��d�H�,�Ӷ�M�18u%�|b_?oE^�۬��jh���o���G)Σ �E~���fT�^��V�M�r�%����ճw�3�<�b��%�'k�j��c�����������;λ��G�n�xƖk.^{�prp�k�1�|������{W��)]6�̝�:?�Wꠤ�)(�w(�;�Q��E*��m@6¨��v�]��w��Z-��L[�����۪�n��݌�������かQߙL;Y%�WN�Ԑ��ǟ0�g�#h�`e*��T'���f���V�7#c�]ܻ[3�n���K�B��Ξ�����'�a�IJ�L����f-=�o��y�r�`�C�`R��\C��ӣ�@�m�/+iv_�H�>�a�Y�9���=�-��C��NI�ժũ�cj�s���Y'<¹�:3�}v��cl?1�	�1�8e��/��Ux+�X�8�(�-敕��и!�������ss�m���z7��^Al!��+Y��^��<�#R�g�+�9��=��W�r����J��A��DBA
�U{%���|@?�g� �b2��
�!�A���%_�����+�z�,�񾔣��Z�[]���;C�_ "G�@�zJ�Ǒ��W�!I���c�� ��{m�z��ا���-K~o���;�|ﳭ��?uw��0.$v��<��E���R¹�J$�1��T���}��w�����a�[O���'�����cf�3洮7���.Ue���4��(ł�4h���������	Z���B���f�.'۟��]y�.Z+�}-��ڂe�I���z���4��~��t��ۢ�������z��d���+��x��ά�+p��GNdw8+?�dD|�j����l��B탸������ߙ�A0�w/�~~2�뿍�K�mҦ����	>�-tz4��]�L Wz�~��S�A���!��S��!�bc�Bg����|g�P���g���ZX}��`�*=��K���� B�9A�O܊G�u9+]	���=K灬F�O�V�ΚK����MM�?-��p5�*�̸֗-3:_���H���q��R���W�=�󁔿������>�Ͳ��281~(+���b}��f�M��Yh쵔� ��.�(&A�g��` �F�����@����"�v86$$�|�<P�՜u������R%8�BV&y� �Ku�<�S�q���<O���׷Ϸp���GC>[�Է;�Q��y�Ӿ!��;zxA��l�OkM���jC&�Uw�U�a"�i	t�߹e�� �m��t��&�Æ�29�T!n�po�u����as����L賛���Ba�_E�1��!`|�;u���C)^y���j �C���}����W�������_�x�PS7��w ����st��%�H��Q�j#4��$/t��T@�Q6�A�"jo�����h��U�p����4�:s0�˻�����	Ҕk]�ij��j���FYL&;9K�l�'5� �˕c����CczW�չ�k��VB����ރYT�sa���{IqI��#�AR+%+�RKQ%�PGc��/�8qE�]I�4B�Zg]��|�ާ���Y�4Sh�\)J� Q����Nmj]�X�8�q�����te�0Ԡ����6m�|�RG������np��E&�	I�3H����~w������E��m&���<���4���c9��&�������~0�m&���o`�	���C]<�Η9�$�nɴ]C�N@iDY�免�HN fE.r_��'�P��O���&�{Y�S��M��Hu���x@���ȗ�m�A]�L�������|�'~�j�ft;�a�<�,���1ɚJf�b��P	D����&��*�
�ߪ^ÁNa7h�h������8������a�M�1_�����ޚ�#D�#u��QJ~��g0�C,���x�5-X�AXf���&se~T���eKW�|KY���i�*K"�8[���"	K�*b�'�6���2�<c"wʼ*��+ʖ�Jwe)��j�(���%lȐWu�b�}D$?/�c�l�	�8#Z|�M�>}�D�"�*jR�Y���Ti�U֏��S+��"Yq��2;��p�-�J�)eVy�I��-���ڢUI	��m"R���u�h|ތ��dC{��\�9���v$�9�[Iǽ�44���u$��̱�qu���S��
����p�544�_(�[MЎ����}ջ��+4���i�����P%���SSS�̄�m	<x�J�I���7�) �&��������뵊u�q���|􅡚�����Jf��kx�~�7�����{Ř�w+D]0E�j�:��hc��wsT#�ʜ�:����C���(���
���f����y�ǯ��|��1�.Q��e�M�{߬2�1��a���Yl4w��V�\�#E�DY��sMy��erR�X�7�܌*��$1�2�p'=.�FL�vC��iHa�˓)���׊q�Ʊ�\^LD�B�����!�^�S�����d�Re8
J�l`����ZU	�4#�Äy���x$R����gq��_f����3gӏ�Xu~��)�:B�A��Q�%C�^�@�$��{��8�����t����F�}}}v:N}y�
�O�:���^���� ���_�"�z*��k�	��p�X���.X��Iw����fr�)t�>�}����}.G�^\��X�A7��Ž�q>�T`BT��r�1&k�9�?��2�]��tQ��ʓ��/���6����u�}���?����~��Њ����I��b�}�`���o�/'���i�,p՗*��ù[�)"���P�S�v��y�}~3'\5D�����ٹn���Z���f�R��Tj����Kz��������X�VE�:Q2߭=�_S`@��C&-�8�yt��ֱ����_>:��_o+ł)_��j�`#%KRq�'�����l?��v�7\�ѡt�L�/�{�<�p:ʷ��m��>����ffJ��FXMû����a�a²�YA��~|���e�^�c���z�����olj:��/��D�}1^���5YͤW#��S�-d�Y���#�
<,t�/?xK[���Y��p�� �D���n�y��x=���u������X�$��~��c���wj�|Wt"��#�������1Y�
���'�Y=My�n���w�s� x�|��7M����T�RX����ef��ks������j��t`�ZU	G�ª�En�)�0�t�m���1P�U�߻'/)2��B�JB�B����?~��`�oY
|�"[郵@�`����q�m���R��V��[P݅}�ÑH��7r&���}�tUG��bb�b�� ;;����	#CH쌟�\ã�w�a��P� ���G�8`�@��!YO��-��1�x���z��-�5��7G��l���Y(G������WHYb�F�;�����y����U�`��#ㆲ[J���e�j;(��VRbT����L��[�:dW�p��]Û>���<+�u��;j�h>Q�؛)��"��s�w�grQr�F�^��캢��~��Cuн^7���Ro�;'#ɪQ�I����S2�=��<�*�uB;fک%\����TthC��Yu�$M 4�ٮ8��m�Κ�S�����`z0��ʃ����l�9�ec~B꺉����u��kɠ��U���)��t>�G��y�v�0C>L+5B����8ݍ�����	�Hi�_��ۈ��z�=�V��`iu���C�}�6|��	H����xV����}�>`3w>ִ�O����|L�T1�>�b��'�P"��˻c�S�A:�c���u���
�i�������f��xr�dݕ���)����*VU����BR9���&y�E�����~�0��+�U�U�:�D,̼Q����ۻ��F��,a�4��������%>i��o��8�7�����VfE$�p\�I��2n��p�	���>.��t}�°��}߻�~C�+��)8뷶U�:���j���ڸZ?����e~{�㿼=/:ρ�_;
#���X�O� \��5RK��1P��M��#FY�Ǝ�8,9�*W�4t/G�pfS'o���#� ]!�3��n���������y��q��yz�˷�H&���_ĕi���@�p�Z5���a��������}�Ֆ˴���GL�5���~D�x�=^�R~���nDMd�"��5�={U�rm������=�uD��v�"0�MtP4��N��d�t���/���p�a��3yG����|��������j�)oj�w%]=�R[7<J��!�zΔ�3�� 7./Q+�/�!���0GA<�w+����)3� dć����܀�D����]��������l�������f�)��x��=
a�Q*�L�v�}ܗ��.��C\���\8�&�!(��������?CD���/����h�Wo��E�ۧǧ�<Ϙ+O�l���2o,iAh��}���O]�����n����x����6(� ��<�w�b�	�|�Ԩ 8^���]a��@q��~����YA��F�D�����m�����F�"t�I��
�x����TJ�^�@�	溯�G�}�ɠ;a����q4��f�2JP�ZyNsx'�^sԿ��7��Ϊ/-c"����d����}�󞭴�b�_�0=��̎���aߵ�a�~��/(�΋�kN�w����n��Ѭ� ڈ[�Aރ�Huckn	�n3W�Y͜���N�Ǽ�Q�����B��v�A������[0��0 ��7[F��s=6����x�,ɢ���7���<�9�H�&,\�!���	��v��z��]�o�m4�T��S�]4Ft���<��l�:�9�)��ĉ�ߕ ���"�9��K�sK����+ٍ�Z�ʻ��-�˴<����YTϧƵ���þ��0�'[�/ĘZ:�I�͑8�iq�1D��p��*�qz}Aռ��F��Xe���܊�#��q˱��6��TB��]"|��k��J��4a�n�?ӳ��~m߷x�k%�TV�L���f	�) �ޟb>u�*����|(%$�(.�ro���vE0�b2�?߾5���9eN���Qv5k@7nO����ד�����c��!tq�;�F�v����f��)�[��;��Ȉ�-S�Z'���(�
���A�S���,���q�ˉc���21ǜ��sPt�<89){i4��E��#Z"Oz;�3Ґr��:o׽�L�3�j(9n���g���t'>�=M��6~��\�~��=�p�������oE�a<�K��$&��X�ٜ����9�����S�$]�
L �d��������G�������<���=
�!hs� {Dvx�DW8��Z����j�Q�ܒ�b�7.baD�,�yI3��t��-�hE�c��,wXM��>קG֤���=ZC?����k�&����? �YA���SX�Ɗh1B�4�������d\F?hjXk]�'��ݎ�7�l����p^Xg�N���t��2��d��ŭ���e�"��(v;�@��y�P�Lu�'��o4ip��d:h�J|�z��v����m�Ρ�s�?v<�Ȱ���̥����h�)y4����߭Nj�M$r�-V��í}���4�����:����1z���"��l��y�w�Prf�e�I�@3��T�U����&=��ݗD�,����{�������10�1&<^�\\��k���+��:���랾>4���L���
8�:M�щ�<^P�����E�=��OCL����4TM,��7C���͔i� ����__�8]3xI����|�3���ߌ@�M�͗Kr-F5�ͺ;��"J^�Bc�U�O�Z�[K=�'P���1��R�:�wyr�] ��
���~%��?O~_�Y��d711���yj%�q��]�$� ڒ�VӦO\�[kh<U�����{T�M�6/�p�(ݵɪT�§�G�+�R^��'�x~O���xv6�������l�����@b��}��Ϯqg�2,��) e�Z��rb�"́c�ġ0*�����|��O�5[lq�𭱄� :��o���s������[���X�մT�&7 �;��p��g��fG�{5Ɯs��˙�,��o+��_��Z��ohm}������^�gW._�,����B�+/�U�Vj�gR��ȑ�EZ�O7�/�r�\A)5�$��ŋ?�cǎ7���)k�/���>�ҫ�����ov>|���ѱ���kmm陛+t\�v�Lz�����uq�Ա���1L{��Z�k�����>v�7��Ձ�{VV��7��~���vz���S�o�Eq6C |�� Zۚk2ɮ�\�X� m���\�k�Z�u�7������kO������w���s�;O�r��X�dW�br�����kR�R*J�: 
�ǌ��fƋ�w�,]��-�~��d��Z��۞���W^ٳ���3_.�J[�R�����j$=/�S�\5ҫF6T���7�o��4�YFa�q�Wz{{���<��/|aˏ.�f����
^~�嶃����>>;;w�Z�8)%���H]������M�g�U_+(��4��T.�=޳��ɭ[�yb͚5��T5��3��_��݇��S��%�x�R{��b�J�dlSK�)%l&I`2M`6�èH�;W�ņ���l������~zK�:����<��%�_x�w����wƲ;�H�E
��ć��V{%� �!jΏ�1�bn��n�����jҍ[9p�@��/���7���b��#p�>���@&W�xV�^FbG���z��Q��Q̾�Os�.B����}�����]�v�VJ`���==��3o���#G������}J�5B�.L}������`����A�"�w��31����u�Ⱦ5k���Ν�|���$���{���}��0�+�������(P� �)�M�r��υr5�$%F}r�X���Z���3���`ǎ��2n�����@z|�ŧ��������:���Xu��r��+$xX�Z$�?{�^E����Ϝ9-�BB�HGEz()
(H�,�X"rEPQl��"6@� HDBoFA�HB��g���9�����߽H	9a��<�	S��{���^�}AW53mJy"M����h�h��N��_I�*�:p��}Ϟm�;w캫� ���ih��14(�IS,�z��B#�����nzP��fp��oj߾���u;5`@f��k�"ͰZ�Ɔ�;w�L>t�Ѐ���^$I6�F���@�CÎ��ư��l1����,w�bK;�٣a�iR�e��2�����Á�I��e[���R��?=P�2e��v��a�A�e@�Ĕ`H� ����B�����E�z^�nJ��ǪUc����zxQg�4.�=�d���!���J )`uhME��h����)π*�PJ��Þ��u�v��q��*ŵ���K�,�ؾu������@K�e=+)cH��'�똱�:s���c�� ۚ5k��G�G33-C^�n\�®]��۶mKߺuk�H$ғ$ɖ�H$5�bѣ�Ar�
lw,g�f��ǒ���.S.��O�j�]�շ�YY�e�yό�Rۖsg�d�vD�&��O�Y�.�i�)���v���Q��bU.��֜W�{��BϞ'㢁T����~����<�s�3jQi�Ӡ<�� G P��"(�(�t3��� K�a�_I�|ݬW�Y	��_�������Ӗ��+7\���_�߀\���c�R%���JzC��x�.��b)�e�DQ�֨Q�Ϻw�~4++�ZgW��X���EXU�aÆ[���o"I����bҮ�_2�h�Q�=v��m&��\��������E�)�$�mѮż��]�l٥ڑ���S��o��*�o/�J�(�34�UD�h!���
<(2r>�@��(r������C��:Q��QU~ˠ_��sfѢ6��Or#YF8b�H�,4E@$�$AG�Ƌ�* �4����0�j�Ҩ�[�3��[A�>qÆk�l�rO���7�^��v�eg1�,&�����L\��(Q�'���rgx��ݴi��{���KVVRtZ�gW��V�K=zԵt�Һ�v���ʲ�H�eoŒ�)�+�&;N2���v̒��D���Ԯ���{}�M��x!	ͮ%�2��ᇒ�Z'��,:h��,�.h�)H��H������/N�u��	����,�~��*,Y����-�x��7:����o�h`�V����n
i��$
�@)@��!��j���7��T��U֬Y��q��ێ�<~[YYY3� RRR�\����f�W�\JQ���	�i���^E� �4IR?�l�jQ�.�߿���~�UpIL��:��z?���HY���W?8+�d�~���^���egLd*&��*���&)jc�V�?8pȁ��~<'����g�e�{kL�ܗ�u�A��i�983�.�<�����d(���<��E�������J���>e�J ��/�T����߶�Y�ԟ�F�\��ܢ<�A� ��� YE^eJ$d��/y\k�:ug����OU�[=~|�{�ʜF۶lWV^֝��4L6�����LÖE�J�uH�0F�L���DLN�5M˧(��f͚/�ӧ��o�=�P���&d]�#�gϞԯ/n�s���lBGY�Ӌ�����D���_t�4�蹣���h�#7�� A?g��\8`@����}�\����f���_�[Ԕ8u�ڜ8X.(��
����`�LVG���,�?*�&pV��)I�5���m���op1�^�c-�~���3�\�؇��?�mϤd2]p��Ѐ�L�Hh�$h@�`8��$DlBa9/lJl�rj�g��o�?^j�u_,�rdA~�MӚ�</��Fc�F\����)c��Y�88����"���_�������-[;ۼ9aj^Z��@e!�Q�e˖e�Z�����3�5Mk��s�'�AE��k̄�h�G������%q'9�[}C��3�:ܜh^���׏<U��׃��"mC���:vF�x�x�h 	F% N�bM.P��>����]��C-O�26jˠ_Fp��3��eN���c޶=ω��$�)J��3�$��j��A���� �������0#㑻~��������][����OJ��SӴ�Q�#cl\8 b;&��`g��P1�j��,�u��gee}ҥK��M�4	T�����E �\�lْ�{��yyy}���hԎel�~1Y�0~L�?�[+�`��������:�jp��[hѢz�¯�2������N#�|�_�E Xb�P��y��6LA%Y�(�Pd@A����Y�g�z�<s������A����g7rs�S�]b���by�{2Ь�(@jȄ
Â�@��@ *EC�� d���_�������UP	��_/�f������>y��p�fZȪ&�ǂ!H�"�A"M+�����O�iZ� ���i;j׮;w��!��o�ު%���[;T&999�9�}�j���R$�1��D����Rz�8q�I,ʴV�X�'�	s*I�\.�Ҟ�o�l����*�{�K/�ٴ{d���*)k��r R4D��ۨ�U	�M�#(F@D�:�Op�lܥ��U�rY��e�/��{R4���^�=w�P��U�2	cи)�(��@Eu 
4�EC�)�x�vh9���w^�R��}������s�C�@����5pp�$&��g��Wp��p;f����8��f2�i���SÆ����cC����V�\������!����/�X�▼���a� >J,?�1�cuC5Ij���:z���q��(�Y]ӿ�ѫ�{={�9T��P�/���߱��Z�<ė��"$��(�Hve�M\4��8� �4����V���}A��Ue��ⰹ�"��z��p߸f~p^�'��"�+�\[p0|$
�3�T,-�`cP�
 ��ry�t Zû�f�n�׭5�Wg�nۼ3�����e���� ���9	�	0���#��bX���
pAT]?����U��u���lu�Ď�vi���C 77׵jժ����'�	���E�f���)������ѰWx��'t]���S�����z�5�Is}��/'���S�Q�P����08Sݠ�ں���D���ZG"Y(R��!��Z���&:v�R�X�eT��-�~��	z����|j׏�x"rτ�J��
6 �4b$������F ǋ�0�V`hG���ft������WT�)77��ݾ��{x�Lޙ�$E�q��fmn4�h�@ <oYU���d9F�J#����4E��n�5-Zп��t�Ҳ�p\�&d���!0o޼Z�V��G��6�`���%{�f�ޑ�� Ef�
�y� 4]ӎ�\��~n�x��;�W�ǻ��Y7eJr���K��#��H�o��S0��q��m���2HQ�>��Hz�~���D�����u� `��� à�|:���?L|�nn�` Nр�T�tC������5 �]
��a��^Tg@�w�n��&�8���嗫�����4Mw�iڍk�˚^H$�@ �a�BD�L�U�p?� J8�;Լy���2�|5p`V��ȼ��:eF ������?���$eEB�������7��5�/` �bTǘ�3�
I���Y�f�G���猌�H~��54�'��} ��G��p#V��m�� ��m֪�$��S�P���i��굙h�*t��v�?��eh��ͻ�Hζ)�H�g"���aAd��a0P�(K2�)��d�@Ui��\;��"�
��a�۲e�G�:=�.��E�+��H� ��gz%��HT5�0�^�DD���26�k�j΀NV7����d�S��-�X������swHR�I�Y��fƘcC�Y�m��T��Z"i�҄X��٠a�YC��բE��8{�{�+�})��׽�%)�(wDn(H8i�Ԝ���懵�R�:�)

u{��-��5k���J>�ӻ��%~[g?��݉����J�{�Ѩ`�5p�<X���!�)*��%)����z�����>��u�f�`7mZ_Ƕ�����`iI������cJF���p�a��쀙/���s8�?6j�ln�>�v��իZT���X��&���ږ-^�����-))��j&�ƶ�B��*�����Q���4 �J�[bjҒ���׭[��`�x����F��C��$��[Ձ#Hp��C��mK����,#�چ�VM_L��դi\�ǰ�%�>��ϛ�ܸ�����u��T`HU]��L"�4��m�|��sɌ�[v�</y��e߽{�wŊ�mٿ�qUպ�,k��6�����
D�!�;�^��ѰS$�FTI9�����S�N����TÆ�K�u*�*��̙3k�|�s��*C|>_S]�MyV�p⋡x�C�ǰ;�c���@��<�c�p�m��~�퇫C�G�SO����dո7)�ԧ%	�<�@�#��tY���� �EB�"�2�}�S￿JpmT���_n�2���-^����-����A^�I%,�$+���,�d��c�E�W�S��F�z��1�}����>͚�K�W�Y12/��H���4M![>ш�U�Ν3�92A����$&�!e�F�}~�-�l�dM�6��� �o��ֳlɒ�;��2��`�N|�����E�������(�>�S�.�!|uXW�~���'HU��nU�KHQp�9�l4���8HРE408�<]vԅ�;�Vc�HKv���e�/�>�D����;~~��;7��ڝ&����d㰮+�ɰ@�P(E�����_g�����3�v�b�1>���w��_����n�))��΃]t��nXk[XXh��+�U���$�(EQ��l��YYY�]{�gڷooq�_��d�">��ɡ7o��h�Ν�#�~4E�
�B��+��1�#_8>�#���P�!�Fw7k���{�oW����>�{�������Kg�Q�/P[�6(� �[4'8ɁNRP�(PP�$&̭����n��l|��+{זA�H�K�����&y熧�L����	@���Uޠ�
@s6�EA:�n�J�۪{����C��1?{��mἏ�o߹c����(�r����ST�4�Xk���ҷ2��Ζ0�+--m��ѣwu�jI/�Y�W'>�䓌U߬���f&u,�}��E'�H���&h�y��H$��M�)jo�ƍ�<��5ՁAq�ر�"�ώ�D��^ SDЀ�I �g�<�$�U�QX���czr�;������̴$�fǰ���w/Z��ơU�K|w�!9Q�u��p~%�u� �Ip�*�'���^����鴐0����Q62��y�=:N'�ZI�X�l6�i��� ����\�ǿ����'x�_޺��s�u��Xff�zZ�ZTK֭[��4{i�'�ݭj���H$��"��Ѩ����x�� �$�K��[��;�Ρþ�|�q�.�{lc�d��?�-�'������N;�Np$QI���BP�'�_nqS�o�Ν�h�n�5Nˠ_��ڐ�k��mgύI��i^�)\5#&�Yߘٮ@�< A���2�>k����+� �~��˖eߙ��hMU� E���4Q�� ~А�!3,���8��,�$7��k��߿����_q:�|u�a��@ގ�ǫ�7�ݗ�HYii��j`ī°�:x��+_0D�I��h;AS��ۇ��u���%�����WN�z:M�EM�;� �� ))	x�P�u�4�rۤ�s��u�FXKy��^-�~�P�������<&����"C/)�� ła��ڐ�렑hv�>#5铴n�>�R��_|�Q���nz���h����h�q���q]Lbk��9h@��}�]�77o��C�ڡC�+�`w��:�B��!��������u�,ɷ�����,X����ј{<�w���(GǠ c��AC^��.�s�0G7o��(Lr�z'^�Ґ@p
`��`�y�"T�� =.9��ζͦջ�}W���م-��7_�q����e_���S�y��^Z.�E1T�%x�B�@�@�"�

��M���az�sk\�0��Y�mݲiR(�G����0̇�u4�h̑�
��董� YR�É��Kڵk3o�ĉ�J1�o�zkw�F ;;�旋�G��4��C~4�詣kl���t�(��� W���1�����o�
���l����C��x���"����D����yaEP� ��@�'�����Mz�~�;p��4y��2��R�.������Y�{�XS�[	X�M��s����*P:�� a0�r��A    IDAT�pP����F���y�V>7;*F����-������p��v�p01u�50���3�AC��w�0C������aC��۷o�߀���B�B��C`�ʕ�+V��z����h���,͙%�hȱ��d��r�F�����t 	}wm��^z�����y+�g�N�aنѵ)�a���!� �! )%8�75.(��rU�Ϝ)繷�������k�����w�y�+��y%U#:e�(x)4˃$k@���!�?Q,2����a�����^�RP�O|��m��Y�?ЍeY�<�+��`0��w�a�����$x=SR��;v�ϭ,���J�]-�o�]n��w������HzN�y�5'�����M�;֪c�L��Mӛ7i��ȑ��7���6�������2����Қ����h��Dp$8ARdPI$��b~7�?ߴw�o-!��ܻ,�~��O��4;�aۛ��@�A1�������ZR ��@aY�F�!�Pj��۱�۾͔���t�����'̙�n���ώG"7�,Ϙ�9͙ei�|�R��ހ9���H�\ѤI�w�O�~� �<!�v��8� �x���֭:}S$�U�� �3�$�A�e�l����(�p[kf�|��;��������~�Z�>��$�4���N��I�k�dhF��((����k59�eۍV�����,�~0/{A��뷾�(rD4��J �E�	 #�M��@($c�X�ܱ�Y�ت�k����<.qIwٵkWʂ�>|�����oI�$�01Cn���^�m+I1^v �h�>�r��޽{��C\қ�Nf!`!�/̙3�֚U���n��,S(���v4�MC�24캮VL�e��w6i���>}n��9�˺���q�tBbX�j�4щˀ�$OBb�D��6�*���G�J�m_�j�nB��n;d5���e��K�(Y�4����?'�qFT�]Hp8!��WHU7=[��2M��M8}FW�v���&��S�5��~�4-;{�肳��Y�oB�90�'�^ Ơ1��&���c��2�kZZ�'�^2`� ���1,*�E�V�X�|ɐ�ӧF��<��L1ǘ��a���3iC��p���$�x����㮵�J씗�Cز�Ӯ��)��q�i.��mgbu�<�BD�W�R�V�Oj���صO~%�����e���+;��������Sg�G{�j�C�����aYESMB��NpC�,��:�i��L~�pe���K?O_�d�X�o�P���6)���ŎR�f]9K��گ�Zn�:�g�~���gff�W�}[׳�����NZ�rM�Ǐ=@ њ$Iz�$�k���"������q�]�������y���Kڴ��~�����i�WCS$㩄��У`��K]��� dp�"�2�3^h0��r��E:���ˠ�#I�޽�C+Vܭ�q��ݨE��f9�i
�a	�13đ�X�(Q�Ҩ��=U�ִ��x���>�佌��m|$W%�bS�7����7��JL�;���Eh�7k����n��`��WN �jЭg���.�5gќ�����1�bnP5�YQ�n
!���,��=55�����\�����)I�}��x��WϘ�Z�{��u�PT�� ����F���pC08�A��2�ޒܩ͓�w����r�ˠ��a��	��\�/��iɊф(+ϙ,p�3H�5� �
�P��.��-|z���O�_ٍ,{޼ZKW�d4��� ��8�`ކi�Up��exs� ����4I+Z�n���ɓ+=�P�Y׳��>|��5kV��|JS�LEQ=�_����1����X��t:����D*c���=j��K�5¶`�c��ؙ�$�툄� D� EA�U�t�	JI�;�/��6�fէ�K������?�~�K`�o�p��m�n�����r=\�"hP9J)V-e��Tj�mG�[V���X�e��O���!�,�:�ns ��!��u�K�Y>A��6��=:�?v��3U}����B�jB`	�������￉e�d�y�5�X���\f���9�����hM�s��ƌy0.=��99�w}yS�/<����I�岃�� �f@
B��z/7��o!a1W��=,����y��mX������K�,������f�U�(('(`�_�	���븠�Y�f�|���-;�	GuR���B�ha��M�5����Q\E��#			��tS�'w�y���~5Y
�Y���{���={��A<ϧ!W֧�AǨ[rr���Z;�o�PUU��;D�I���a���g>���g�g��S�����k;l�6�6�@�P4� !�}٬��~xgܼ��|��A�'��V��y��'Pg�G;%ٙ�I) ��9�5s�<��Ca�^h�/l�3k����e��5���7~?AU�V�瓑B2F%���8&�Up�Ǵ�y���nw�'�{߲p�+��2�-�����/�X;''�qUUo#I��ٯe�L��I{lM�5��Ғ�D�t]�GR����'|Ӿ}�J'�����/��qt��I5u�v�W��R$��!�ۓ �`Y7@R�3t��/�խ�Ԍ�C�H# X��h��������O<X��k� �$$A -�G
T��0MC�'N�۸��۾���{K/�!����ygF�u��M4t�f����C��)��!����7�����2��.��gQt�=h��k���_�D7���}-,b����7o~���0#�n����*4x�^�x��c�$F�a��))9��1cZ���_�{�u���3R4��=dl�
"ρ�� ��0��A� �Y�}<�q����^K������n,�������{�~3�:S0�>[X�C�`c)�(�ʚ� �M�&�i5|.ⴭ7����q�J3w�uׯ]�LYY�`�ݞH1l,ck�IJJJ��Ѡ���6!B�����Է����R�����7�y���+W>����$k��:�r�Q�(:�JK��������N}��[�7o�l���`�:q���I��'�_s����E>X�`&
!E� �@9C~ok��Z�<�'�x�n�7�(^���v+ܴ{z�b\o���5�,���F��AC�A�y(���Bٙز��V�xj�e{3�����V��֮��j� Y��0��p6Ӏ�Ipf���3�@XcgFF�k��z��Lk[��˺���%C��w߭�nݺ����FSU�9���$cN�N���&
�����R4��A���_~�ͭ�F�;gNگ�s�J�G�#r"�f�Yh�w��T\K'	\Y	�ͯݱë⭷^Մ3W�A?�x�5G�o~=9��"�K)���%A�e�#QiH������f�_�Z5��p{�啙�>g��Z���4�W滍��d���4et��c�Ɵ��Q�� ��o���[o����;F.��b��B�B���9sfʦM��H�tO ��!wU�M�1a�W�vhZL
 �Q)�}�֭&�cګq�)�zҔ��_�&��zxt�u2$ФN� 	N�9�!�F� �����]�7��oq�uW�A/Y�9�U+_
K;eE��� A�� ��@r��<��Pj��:��VjF;�ƬY�v�mRTJ�`�bX4̀P4b��1�Ԯ Pde�5�Z�t�w썷�[����-�4�~WU�h��:ao���ںۉ�j�����0b�(X���/<>a��8yL�6�v�~�����wvZB8��Bi5<G���4C�6J0�:%��J9�[�U�����҉��
�W�A����ݷ��G��cc�"�U5tB�P(`*��涳�s"�x���a�8������sK��^`��y5�۴���gΎ""�.:��3)�$��#�d2����Qn���-^�ѣ�/���q��\Y[ױ�'f̘��cǎ���G�4W�$i0��<@JJ�~�q̬t!�/+�>�n�:f�#���Y�,[����e����\iy��!�a���� �8�
n�I����]EG��FnzǑ�uU��^���~Z�l@��ѩ��@c����,���!k�� �%����-�l�b�G�.���`�����7=TPX0�e�t��S$mvV�KUԘ�
x�d�
7�i��ŗf��G`���,,�h�srrVemt$"�c��,O�I3��]�"��ܔg(fivqϛ��6z��JM�X�7N}�y��]���jOG4��Z:!�	$��f�Mr��4(���1Mꏯ=��M�7p�8��W�A?8��Nl��zBH��Q�4 0	�,���@�($>�(�;�k�zi�w�2�ȥ �|α}ݺ���?�����^�fMC.˱:s�HQ�d�µ�H$�#	�����N�6mZܭ��&�>�� f�/_��xQ�������Țc�s���*�8�����仼�/���-��R�J��������Qg�NJ���6C�UP`
ܢD�xHH.G��%y;�{��ȑ'/���z�Ug��}�����nx�=S<0A#Y�1B3@�d ���G�r@���o�ps�J����999��-������i[3�Ή��p(�4g��yEQ��l���5Ͽ�j�%��k���B�J#0}��:��o|F�ۊ���v�`���S��ib�Q��q�(��N�������|ڶm�J�6^,N��]�r`��'�C�QUNeI�?Kْ܉&�'-���E4�R릿Ԩg�⫍��2��ۓ��X:N=��[�=6Y�h  �4�*P:	��C�堄�&��o��I�Tκ��}�ď?|��Ǟ�u�A��gN�P$��QYK�145�*�֦�4{��_�m��/v谎��/{���~�eMQY���*m("�"MHƂɲ�$�g�;D��u՛q�=c�nҤI��],�9ϾԺ 7wF��wu(*g� h��do"����H�<��]l�h\���jӯ�n>�X�tPq��/8%�Һ��� �f�!i`(�,M���)�sQ�]^K=��b�����C��|�e�Ν/�lBY�I���n�"k����0����$!j�)ޤ����}����\���B�B�z!��\w���)�$w�eY��8�&L%W����dY�$%��}�v&O��#^�������o��(-*1m���I\N�)T#:��KUiJ����}�|�-o]��M$�b[�UcЏ.������g��Z'.�!)RU�U �dX��WⱭs�j��k�=��ł|�ǿ2uj�m���@�"(��P;�rfIT,��HS�\�I"�Q�F/2h�Ug~�([�YT?���żJ
K��|�$F�0�Kڼ�	fu�/b- �"Rhݐ[o}vԨ{*m��X�}�q���6LI*��F57��`Y\"���y���N 	X.ղ��~x��^7^��*z~��:��Z����dP�
����.B$���@j�),/����tӆotu�r�aC��_���>��r��)���4͎|�f�(��C�A�j�n�X�fƌG��y��W=���~?��-�:۶ms���[���S��4G?h�%9�����zM�tt]/!i"�޻���W՟����;���x����ґ��;`p%��Ns@��dd��Ϸ��7�)�%���&	�b�C�7��﹉{,�����UK�^�&@�d3l�J*$#¹H %�W��1����zzW�Z�'ｗ��֜g���o7H"�p\�B9T�?hβ5#Vg����R�N�iw��xTT��kk!`!�#�z���O?��޲��{t]���9�j�26�c��JK�1�w*!!a��O>�q�ƍ��ۣ�ٮ-����T�ז�:d�8'n��a�b2�(14��HZ��MYC������jmЍ�\f��-}|{y���:4@ULÈ:�j'tn/�Cl��������Z�J�]�nY�E�>�wjM1����H�2;bT����cf�j�r�煏F�?���],մi��1��y���\�d�S�px��iIb�1C�h��SG��ِ��f��X�~��/���� �"��)��������=�F;GA������@fi���E�_9�o�lʭ#�U����V���6?�q�[lqy�d�"8EC���p�ˊi eI����2��x����nx���wWʋ���u����!�|� �>n��L��L�p$�Ĕ� ���I���w��f��ի��7N��,,.�7�|���U��Q�W�$3�C����?�Ǚ��R(--�����o{��;��=�ٕ+m[�"�=�B¨�S��.8��M�$x|���T$)eJ�����|y���Ж-i����(���)��) @jP�!)@S, �B�$Eq[;}V�~=WF��a�ĉOu;�����u� gjs<2�A85;��.�i:��إ���{yԨQW��Ѕq�QW�=�ص|�0�.�p���t���gRR��������^^�+NNN�?l؈����{:������'7l|���tY���cy/rv��M�)� E��J\#\�xB�w��v��X-:R���|Q�����V��D$���FT=�Is@�v(��ߋm�{�0�۷��B��;ǽ���M֮]7�4����0=q���P;t��A;(%Iju�޽�1v���:־W'��O���ȑ#��i�5:8ƠÐ��l��q������~�N��/>�̤%5j�0�ڪ�f���+.�);�rYi�@�&�-��z�^��� .���D�����h���­�[�4���kS���|��'�D	�F�=¤KE1��%��(('�SA�my�.S�G���z�K?O�⋅υC�a,Ÿ�aa�=ΜC�H��dLϜ��$I���������?�Z�����g���lذ�;s��{"��X�����������r���ɷ���[�v�>n���q1���Y����S�ۅP���$�������G
I
 &=��o��{��v!m������۲�N�n�!;1D T%S ��  Y@��E�{g�F�:Oy�R�v�����÷�9{6�1��jb���ֳ�c����P�<�h���]���aÆY�1�­c,�r�Ν��v��	>�o8A^��1
���S�DBf���s����I��핬��qQʶb�ә���t�B���g�P���$�Ϩ���O�Ci����c�e˲��,��A7Ν�o{��ڱ�ϻ��vU�0T@�E���� @	{�����u�
"3C.떛��|:����N} �a,C���P�B�1G��$�x��oN�0aa<Q4^V��[X�m&O��|˖-3H��A�4�^:F�V:--�v&Ǚ�xUU��\��^ziƼx��.\�x${�İ2���v����$���o��!�qp��rR�\�dҰa?�m���je�/X���m��4����4���i�n���à�6��'�P�]�玹}��Vƻ�6�����VYiYoAH\p�<��.,,4׳*��X�;a��>5jԇ}���j�+�=Xװ��@g�w��:s��TM���z:z���*���X�tA����vO��L\����x{~��	�坓hhR�ƀ�.�q@RD)BN�8�q��xH��D�2�Wf[�6=�aC��k�y��0�����(�5tC�t� HZ ���NR����N�8v�� <;;;u�W�'�+<wǳN��aΆi�7״b3c�\�1�\T��=z�C�T��Yװ������믿>�0��t]O7%�%�t$�p;�1��K0�+��OF��V�>�V����ٞ}V>V������mФj>/ڀl&�{� ���&t��xҠ�?V�7^-�aD�9����Sh� PV� 0͔D%B:H���TKx��q��nzmzNe:t��ګ/�>u*oD:
	T��E#����⺖���ɲ��K�.��~��խ�Y�c!`!p�x뭷�[�n*�0������b��� '�(�,���p�`�zO<|]f%IG_2+y�:�����������!�˗�L�h��!����E���׮:bѰa�T5]�s��c��A�c��N~��W@�
J�ZIIP*�I��L��k    IDAT�ぅ�j@I��z>n7r����+�im�����ضk&ES�:P�,E3=r�jǙ2���$� �ۛ6m:��7���w^���������� 0v��.|�a�k���q1i8V�ƛ�Q��&�ʑ=3o���#�?�s_�}�K?��q��D5XC���g�xDt ��ϑkk��1�9`��+yϗ��qo���9�;��~�Q*�oiI��G� Q���9یJ
�D�������ӳ����R���?�<}ɗ��I�:��(�Px�f�WaF{$*��ݝ��w�{b��{�wq�Ν�F��R7J�|�����k��6�0�{���c��H��� n�3��KQPPP ,G��X��#F֧�r�.��W�3��:��[�t� A �� o��h��y�Qcb�{.�N�qm�1Ծ���~���G��Q<��P��>�C )2DT��C6>�nR���޸�2�������1�Ϝy� �f�K�5g�83 +�,`��!�3���y}Ĉ����j�X�����ٳ�-_�|�a7�n״Xֻ�!�,r�x�v��*�-�y���fT���O�d'���'�uu�=��
		v\"�@#� Q��$%�aԼ��?l={VJUe4ɸ6�G���֑ի^r����!�ua�������tā���C@�NB������Q�A�*�)hܸq�~����I�C�	oXs^VV���v�q+�rԆ�������F��2�u�˃��q����34M�C�Ã\���c����E9ES��6x���w��<ws����C�{�Ǐ����1a<<�^��q $м�Y�H���>x��Kw�+{��5�ƾ}⺯�.���_Z�� Y��Ȋ�o� !uj8*A1�'�P$ѽ,����v��h��Ϛ�z���7�"G���a�v���c����!w���a�� ~@���C��IS'N|zi�@���6y��� �Ƚ��������%#��I�h�1���騣A�D֨Ysܐ!�7V�����O>�ꛩ5$e�+j�H�
�N�Dh��ˀ�r�����|�h۶Z�ǭA?�ه͏n���'�vdX� ��!"�A�� (@A��!b���z��ۯbV�~��3��gϞ�P$~�0�dL:A��� Hp���s�H�Y�4��������z���f��[X�3�ޘ�h��կ��'�����ML0EN�>C�%][޾}��'N�5�}S�a���z�������`�5Y^
�nD� M�hw��� <��6�E�q��<X-J��Ҡ����4g�|A�LDM`TD�M�AV�uªa��ÝU��E]~5mh��L��T��;w�+�lm0��TQ�Y�}���@�u���1l�w�Q)���$�q����z��/�O����qlMW 556�L�-.>���gH��1��;?�СrD�.�W�I/޹{zRY�P1b<<� ����p��$ǀ�5
����׹��ωV�Bz��r\\��ѱxӮ��:y-g�@�*�<�`4E����Dј�.���_�L�IO�\���|n�҅_��d} M�6 �б��ా;���T��׵���oͨ��x~����իSg�7{2� p���j2�\.��3��1#lnݲ�i����*?幜{�'_��睙���i6Ё137 ��+����4=�-�t�����OU�g:�{�;�^�m}�-�LM�n�K���p�*�$A�4II7 D�PƳ�ɺ5��~�m�33����쓛����7��|�A#���u�itM3L�d\�¿�x����~o��qv�СZ�\�ֱ���O<�����3���t�m."�u�e����KH��}۰�\��{nZ�����R���J$���r9@D���@�DI���a�A�i�� 2��G��]1��a���9r��TŨ�aRM�hS%T�� �4�Qd����ݤ_�i�G�����I�����?���|{y ����� ��Er%˘p�crŰA�&�1f�j�t�9�τ��ð�^�D")IIQ� LA6�ho�o,�9����&YUEn߾��@XP�����{��1��　�$��ԨQx�5�KR�}II��g}���J�ɿy���߹~\2����1����N�h���.�9��2��%:����k�=33����ʠ]����ks^u�B7�0)Ҕ����o �g&E5S4�E~��u�Go�1�R��+V,�1g�'/�1TS�cx��������g�5h���l�O�Z���[�m��m�ڽ ���k+..�KK�����B|0�sCa���rTJ��Q�UD�&YC����tu��N�FP�BӤL�T��(?M�E��	Wβ�/!��ټ���U���d �V�,�j����>��z�.�AQd?MWxtDp�2)a���P(�)z~���^u��U��}�3�ە������QT�q0	n�l� ,+��$��c�C7��X������qōA�2�5����,	<n�289
<M�Bf\�<�
Â���u�p�;�{�\�ޕ��'L�2�μSyϒ$]3�S���:x�v�X7�����RRR?9j�x`^���U��o۶�q��1�?��gΜ��B���j��
`x���UTգir���.0@ ��u�6�B�GCG��^���@K`iH�b`�A�߉�B�$�(�0!���(�*%��Qb�9��θ\�����B�;�W�fM)!!Aʬ�%�������0;|ܸq�:�"a@lghf�Y�0aάM/*��z������[b�Pl{Ur;����}^����<�!�T`)���8�!��[<W�qN��ց��99.n���7����s<�P�$�ZS�&jQ�4��������lJϼa|�OV
O�+�Lm�)g�,� �c6;6z����Рc�	~x��~mf�O?��'�d�n�X��s�g�w��e���n��5MKWd9M�4������a,�c:�A(�
���:`q��"C@�?��?��4��4̀�,E@�?	�4�@��$�j �BS�JӴL��d���H�*`Y�`~w��\ޔ����&M���f��\���9s��(�)+Q�?��0��tT�Ͳٝ�v�2nܸ*�Lf���}aXZix�3n@)Q�Q$�x�6�DA��7��_z�o��w���x}�qa����w�]��<��B^7M��&	�dUU��� ��������b�y�˞�u�ք�^}i�nwK������`�f�G̙-wQjӮ�㯼�ʶʨ���FO��n�|�رB���|��s��E��檪��u��a�TUMTŦ���asL��H��C `&L�z%a� �4ɀ�+`h $M Ks�&^St���#f�MV/U�A�U�J�$�� ����.������+��i�
�2M���i�-�(*�$ȓ<�t�~�x\�������;v숴��v 0u��v��1K��X5T�$��q(G�m	�(�:�j����{_v߾}q�X%�}�έ{r��َ@���4(AW��P�@0,0.7iʜ��J�:7~���]
��~x�Gm�X�i�W����u��l��ʃ�G$ Y�U=�zV\{۠I�G��Y�)���ٳ�0��f�v�2E�L�W�b ���/p�]_�3�WP\%[�uS�����ż�C�g�RԈ|C(hG@:A�.E��h4�+HGe�o��*�c��n�6Ya�c|1�L�����c�U�h�0��D3�ɘC'@Q%�1J�f;ğ�K���Mw߈)�iN�����(���$fY��a����E�����\�\�f��C�����z�N��u��%�ᇓE�C�dwE]::&H�������e��w��y��?~���%8)��m���xGi�X�$�
Jy�<��/��pP.re���ׯ���y��Kp�J?E�7�Ǝ����O����������	���=|��꽧{f�P@���'j�&JԄ�!**���l� �����@�E���FqI�*n��20{�U�U�wn��T�'��a�&�~�yz���]��y���-�\N�`�9���D],!r�O$}�E�.�w�E�)m��]�|y����t����^��I�L�)�b��9ݮ7N?�̫G����6_����x����}�YxÆ/;mپ����������-�L���߰Hk-�7 �\0 m�8,8���\4 X �<Z7�^�*2i��� n�5�n�Chi]j� z� ���^��6�@	������ 3+�Gp	�Z��/�ݡ8գ&�^o�����\�k���AII�[ݺu�r��6��߿�T����*�
�M����+W�s:��`_�~�{�㠩�>�¢8Ŧ@��ȑ��<����t������'�	Q��	�K���0\.���D,���^�K�'=����t��'s�����,.��#Uh�.K��j���BSѐф�zw�ŏv�\п�O+[�~�g��im�f�-~��K,��ntC�y<�l�=��]E��9�G����o���V�l�p�ߢE��_~����o7�O$�Sq�PD�L*�'��Su ��	�|�ˬ���/�p�ɝ�$��0���� ����Q#��Kj����|�v��&�@ ����-,�z4--5w��?�T$k���w|�v�G���TU�;�N�ñ��p������^��o<���{ ����_0�ׯO�0�d29\U�
-m�����;>�2I��t=w�G�?~���:��K���]�����P<)q9�G1��$$T�G��͆�b�#���Vy���,U�U�u<��_�o�}w��j�)6Dȕ��#}������"�cH�H�Cu{��o�������cŲ����Γ�p�E��Yݐ�sh�0����[U_��y�5hР6q�m7a��wٲe��k�)ްa��D�$�4�f� -���R� ��Z��_8��5ov|G0��.@�14���N@E� S�<��u1�H�ڗ���@ �g��)P��r8@�7��3d;��	���o������ק6es�M>��C���zEE��#�<���/l(�5m����y����+�ܕ�fO���{�=�;^M�Fa��;!�)�~���N+����ʕ��/���;�ǧvH�=&|NS8.DP
W�HԸ��3�Y���'�Rz�m��䇯̿���}���G֬z�
={�O���-�.S$3i	�M��ȸݢ�0����Eg]q��h�|�|�Ad��ۯޱs�G�Q��4)�����$4��hV�䘾}��6cګm!h�Λ���Gy$��;oT����ӳZ?]�7��L��L&c%�Ͽ � ��byH�ߵؼ9��:��w�kq�8��(?�S�,�n�#e��C;B�C���d7��`R����w�����)��vS��m�=�@'У����C�� O߅��04;�NĽ�(���hɋ�z�7�^{���l�k/���N�8q�;F�<�J�k� �`�CS������|��u�m����O�w���W��c��é����p�p8$<�C�ለ{=b��z'���Q�/�t��I/X@�v�zŊ�}[w'�Q/��.��h�ń�P5Mq��h�xV�������h���g�8���}������78��Т�~6��Uq8j:u�����o�ׯ���|{��vy����ﾻn��ƺ�u=wB.�=<��J4M �h����y �V�0h��hV�ٜZ3A��E��Ej�O\�ݩZ&�.���>�3����;Im.7�m�  `����Ҝo"����wyv{�����}�gNI�3���md�RP����L�%�E��8Y�T�N�FUU���<�>=�о5�̂�?o���s������_�����H��.I�B����4������n�k�i�3��੧��T�S��3�D�Z�����eѴ^�5��v���/|�%|E�"�UECȷ5ѭ��'�����^���f޼#7�����z���9&�}^�4��tр�E�jY�
������U�\pw�SZ?��_��3�����x���(BF8��/�F�IǶZ�'��z<o�~�i#F���o���>͛7�d͚u���L&�)�����T*��d����-��J0d4˜ �ߑT�7�S��1l�Y,��l\��!R��;M�vs=�k _#oz��M�Z5}�$�Q�`bZ�>[ NM�������?���W�:��YK$D<��@�?���p�\M~��i��z�Ӈ��o���������]O�2����v�4�yU���p��~����3����}�1�n���
u������-u�+ҹ#�tRx�B��Q��E��D��D��ma���c�Xrƹ{Uj�t0�_}��Qj]�5��r�5�z�b��9��LFĲ�hRݢ&T�Z�c�sք���M4nܸ�׬�����9fP��--F&\���f���6t(-�7n�z�A<|[������s�����X�Y�D�繜�SӴ�L&��:<- UD8>��E㕇: �� l�y[~n\k���2C��(#M�y &��!Ip$����	�$��Is��P6�R؊iϓ��X3�Lx�'�>���_�P����!<V��µ���Y���$Ǎ�^j�i+�!yA�?���������áG���u@g�o��w�8/^��G�ΊD�g�R)�Y��A؋�{���QSlc��#�	'd��Kw��e��7�w��~L���"S�E�RhuB"�����Cρ�]]6x���5�mQOA����Y����y��G�٬�"$�0���2,���Q������b��8g��s;�ҷ�S����Ke�Θw�ajZ6����l�[�n�~%�0�H�s�:��ACډpmq#�J˖���ʇ]�����aB��f��\.���nj�<\�� �����vK턚7A����� J\�xt�H4#�Sӧ?���o����4r��HY��,���]���=v�� ��z@y��dɐϤ�p�LJ�!�}P�ޘ��ə�;�@���?��뮻�գQv�h/��g )a�6�܍�6ߞ�f������my��$IM��a�t�O���PXz��Ǉ�[���JBE8s�()��g�
3��>YY<c�N�_ٯOA��٪��}}��{o(i������� "c�X��u��ht�F}����_�Q�'���-�믿��{�}p���=��4��AZB�ׄ�Ƞ�8���{��9n���nbl����m�\����3�Tnݺ�d�4�'ɣc�X���p#�2[�d p��-���tK���2 8��	�����=��j�,r�����>��8Q� ���o�0$��7��) P�F]k��)�P��3��� ZP��	� ���\��Bȉ55I��+J �%�p86�W}>��N:i��_�W&���wv��ࡇ��'��4L����*��s>�u���,R�VS�3&O���W�^��/>�������%���lFx�!J#Er<n�_�%Q��ru!�򲪓�/9�&l���G9h��/,.�h}=��u"�Sx��54�XCJh>�h�'J#��v�����v�r���7M��t���� ��r�D�N�CX���B��3�;�҉�[�'��v��Z���.���O���7�o�扱X�iXZ ����"6�c�� E?25m�i�Z4�b;���8;H����� gşԩQc�DY0M�z�� boߣ�I!�&}|G����������X}��sf7�K��bխ�-���w��!v��Y�G�!�N��k���������3�l���t����swv۶_�����}{�nU�k���A��C����\<Ḫ�^?��K��Y����ڽ���`2���(����p���P"�A�hx�d{t��%��׶���[+(@7�����E�M��T�j"뱘�.]��hjL
=�[}�[���p��7����ׯ����O������y���Z��餕�ҩ��=�?��kgΙٞ�}קw��Dz��_}�����dҙ_�ҙ��x<H�4���C'�<{g�&ӝ�5�9�W�i�ri�g�]?��    IDAT� ��v���۳'��ٝ}E�l��<�FS;��vB��������Mз����?�qg���:�iZw��F�Gmf䘱����D*)5x�����@�W�(⯑H䑣�:��v3�nv[�<�@�gW<;ӡ(�!G����.�� �1X[�4�x��[��n�#}���2l��`_�{������e�t�/��@Ȳ�y]BErQX��-u%�[z����-l�����-����%ӧ�r"l��6��Z���sS�E��Q_�/�?�;*��Z=/����(����sF�T2�̲~�1Ǜ�������|�]s�Ig�A<|=#Օ�����_���'.BQ[[����K�36��B��/�Z��w@���r�� �$��c��=@Z5]1�;'�c����۵|j�v_%�� I�5�{���ќO���� M��pX΁���&�!A��~
v!�D@��Êm�����W|��uI�jlnjq1`,8(FQ�d(�l��N��,9����WU�}Y�
�!h���u�����~���C�PW��x���O'y��I��p�?�;�j̈#
�T�׌���}9�k�8�O��> �a�pB�"�sgB�;�������ւts�:��'������SÚ��'�Z�D�a�&��q��LazCb����r���$�̘�?������d2��k�23-�ycLjMxE"�5�~��3f�����*���V���o�޸q�EF6wZ:��i�4�#�4 $)�)z�Y|��?s4C�F9�O%0|Q�ٓ� �!4�-���`'��������ۉq���&y�C��5߷P�gY���;`�?�B��S����Z��J�b�fV�>w�)�٥��9A��s�H����d���w���7�[]x챇�5fL������f`�ҥ�[�t���.�˅�Ǻv(+���� g�߄��ƞ���OP
��w�>�y���4mߤvA$�q�p��"\.X�|>��������=��Ў�^���Z�ޛ���/�\���es:��s���)t+<H�"ψ\:'29��r�%K�O�|�e��O9��Y�8y��gMӳ��\.�8dl>��%m4Ƥ���<z��1�����{��Ֆ}��������NO&��~H:�c}h2�#yқ_j�؄�Ѩ�d��W|�XF�pQ�o l"�p�8ޙt�`l[��@?�����,rj�4�?����:>�\K��Z;s�Dodp	px�5
Z<\7ƌw|�C:��I����n��盇P��HW'�R.���0|덍��{F ������:�g��;><p����������=>6l�V�|����kƪ��k��	�����%&��%|^�#pk���o���^�~啢7�{pHe]Ӎ��(v�3Bu("5��PX�PH48]ۛ:��y֯�Tz�.��

��:}�qM�0��tjIa�Y�yD.������0Uw��N�gmѡ�9{��E��bZ�5n��c?����D�`lp t���)V ��p8LU�����㯞:��M��[q�{U�8mŊ�n۲�R�4N�oh���TdJ�n+���oi�X7�	1�$�A���D���GfX��:|'�b��o����&0�Nj���ɛ�i�G_��OӺ��F9c��/�I_��Cۨɣ>��!uԨ���-�����xi>��$��>�+�С��+�.�<�֡/�<ic�|y���\�(j�օ��0o�x�ؾ}���9���0_�C�8��.������/������{��g�:�i�i:�d��Il���L�$�d*�a׮ݮ�;�ނ��~��N}��]�u=�q��.#CDJ"2�R�69��F�s��~3'ܷ�C���ۦ  �������|;�F8��@����N��L����EL�ѭ6Մ���<��ɽ��ou�Y�N�<)k�t��Hj����R�g���(���k�N?�{�9��鍴'�_�pV�U=u����r�q��i��HK��y-��Ֆ�؊�ff+���BL )��0��������C�@���� �Tcj����;�BG�5�6��*F���Ȇױ-j��O�q�\ΰ7�j'Y�ccb
4�c| tFP���ʆ��� ��$�1�F	���3r�oma�I��
FSQQ䓌�Yԯ_Ջ&L�+��{�Yh�6�~�m����zǎ�Q^�].�Vya�ce�\צ�Q[[[W٩�����;��s�i�<!?t^�qW����1�<��
i9�W��8E(�!@����� ��=UG��zր?���._����s���,*3ǘ������p�BO��Ҭ�x,-�K4�=�=��x�Eo��y�SfT��Օ��.��.�[�▱9'V�K]��z�zT�>�i��_mo�����oϯ��yaV����L/cc< !h��Хؕ�:���o�?@Q�e8��ƉȄ�f�y�f`c656����9����!jQ֏w�é��4�p4{�WZd,m���f�HG�؈�=��IC���Dv>�|h_���Q_�<�A+?|�HY�]�_��>�ذN�ŎG �c�`���A�f��.�;oN$˺�������ڳ����~�̙�z��{���S�+nՊ���(�,0�M�L�̭�_�k�Μ�&�B~�̬�ӟ:�yߢ�*��y��D8��E$�Tު�����sY���0?����#F�~�Կ'��q@7׬����+�wN�Na
=�	o�/R�0�2�1�i_����z�Ͼ��A�Z�X�5k�M�1e\*����p9+�'4t�n�[���r׆�B�^5��ڙ�C;xlɢC�����d"�s-��Դ�Br�? 9��_�a��qZ�▯Y�����)U0�� d���p/�K�p
7j�Ԇf ���j�����u��`L?6���}�A�L@�x�< �d�K�8o5���L0'��=�L�����^н@K��Q�Zy�� -��Q��1��Ң �����_h}���M�-\ ���\5���N��Y���f͙g�Yp�P��N�gΘy}�)6�0� :�h�H�-�}��<b�T�:eȐUUU�gB�6x��u�Ŏ-[&D�}�٬y]"�u��@P(^�P�Ţ>�i����I�S�W=����〾�Ǻ~��s�bz_:+|��1���gc�H���}/	�\u��=z��F��k�̩���K�w��GcCq��y_�E���.�p>�{�9���s�,H?Q+NQ�W��?�)��C�������4�'�T*�OӰR���N,�)[����s�8��Z'�Z9���	� (0a����������K
��� ���$��c�I޳��i���Np��ng����⨇�=�f2�a��9��I��!,� ;����("M�~�u�~���ϵ����M ����|R��w��64�ɾB�_!�����r�).-����7��פ�l�3f̑�>�x�����af��[ �/=�I鹜�~?��#G�������xcڝG|��ʹ]r�	EzVx�����"��	��#��)
�m~���'5�w�Ymv�����ꓒ_|v�/��9�O������dL�(�l}��d���ƞ:v��b?����2m҈���Q�i"E���B���T$;����j�y�O6d�9��b�#�zW/yh޼��W��ն�5Ä0N$~�%:]'�I�m��2����l�NE:C�𙀇w :���OP�ܠ���oL36���M3=���R�� Ԩ=15c�_vင7���Z?� �A����6���O0�;��ӳXAlB_Q�j�<��1G���d�f�� ]�Ⱥ0f��|zh茣��w��tG� �I/�����ɧ�M���?����8~���c�w�!���-[�ᡅNs8�3E.h�+4
��N�y��A�r��e�e#��E�HH�����*_��)]2��%��Q���z\�����O�h�ȄB8��#�~�GV\v�k��ڍ=
�V��|���k��M�{��P���n�[47�Es2%2�CԘ�m�>���ҋ�8�DkO��?���/^��z~J-Gu[f�X���)���|r���g�=�[i�9k���3���ի.�^��R��u@6�u���!��py��$�ݦ�ZHi�<؄�m ��d�[��<s��#���t��ONB�.�k���?" �n%`<���F� A� ��Ч�rԾ�����c�	⬋>j2�i�MS=��}���1<	�� ��! a�b$9*k娇��9��A ��։m���/��:��B�K��a��bm@FdT�8-��}�{���O�8��]p�y��u_u�gm�n�L�=�^���B�>��#׷��V蚖p8�����_�t�W�z�����5k�^�s-;GGSZYD�D@1Dq( T�O(Q���PxgS8tg�SO�[)��w��Ջ��Y��{"���E�-̌.�N�0��0���)C��Aߪ�9��on�s�M�t�s����L���	��������!��lTU�3_|�����o�S��VWWw~�o�\��_��f�e�) -R����r�r󷒓�Z�� E�`AC'��!Nv7�@�gO�]�ZP�L�ǃP����=@`I�<�e�v-��4��t���-�p��i~g����쬟��]��	��7��cl Q�����v�=�y�V��5�����Y�9�CDK��#R��V� U,�}纪�W��m�&x�̉����e���>v�qG-��;���U{��4�����?�xg2?���nFTRR"���D�\7�0��߽�U3��yg75�۪�㸛�j�}~o����.E�ZJD�A�����8*r��0����X����&�N;�`��{�͕+]����9�7gF��.�LNŐ��TZM�I��)"�s�&B��.�d����		/��r��s�G�W�Tʅ0�D�ɍ���^��UU]w�!�G�s�=��oO|����W4v�خ�]s��i��d2��	X˓��3w[��tF�,��P&��M�1I^� @��X�#G��u� �j��r��Js�3��E�fF�D=}��Z���5��κ�n����$��{

$�qO͜�w�	f�!sR3Ο�N��s3ޜ5��@=�/m̜',ʟ��y-++��Gp-���&-�Γ�'���X���m�&�f)�a��n�y����m�9s���V�۫�73�t��_pI]}]�GU;�+8���iZ�ۥν�ڑ�;��B{?|hY��<6�2�9;��%*�"�o0$����7�����_�߅�/ԛb����^*[��S�J⩋BZVu"vե��0E,��qM�s�H������'�d��bo�}Jժ7ޘ��zl4��#7�uA�kll�F��x��tѨAm��o�qZ'����{kFe��o3�\Ӭ�f��X�e	Z -;��ӟ�Xn��d.���rh� e4��0�s��,��ϱY��5����/��hoJ���5>�N�\Ș���V'�3�����S��o�P5����/����͉�wt�M���2�/����U2�1��#ʂ���O ǜ@ �Ə����B��@�,v-1�0���$������p(�bYǊ;,X�q�������<yr�իV-�匓`Y�}��^�*ׯ����z���;�#����B���W��;���;4$&�b]��.T�A�WD����\4*v��/�]+�8t��m�������5w��k˻Y�1+�� �RN�ý)���!�nt��;�'��3��V'�}��g%7�z˭��d�Y�<����p�O>�<ݸYC���+�O�~��nݺ���c�s�ر#����L�ܦXs96|ա�ȭ�e�<�GK�u ��(����%��fh �F�{	jVF9t���<+�@�� )�����(C:�d<2��q8�B��tN	s�u;�S�E�R ͓�(�`��`�|f|>ƅk�\�B
M�$B(�� �Ƹ�d�c� `�Qk�6��C�C?`�G������,�,��A�;,��aq�����v���E���	�����k�[�red���'�c�+T��z9]�|���\#�i�N�wE���7WO}�����_}����{JR�#=�{�zD�?,�p���H����>��YJ�f��#���X^}��3�-[�+Ni�]�T���񤈧3B�)��0��"��g�rY�0.y��z��0�P{���YI+��4CU=o��W5��z��{�SX����}���F
E�m"�(�q�n�ڒ �[�mKC�br�%M ���p�{e�l0 m�u^���Z-���k��t ?~'� Ks<���1�8���[Nb���Ǳ3����C_:�����|ƍ3��ˣ_����Z2��"�ӺA� ��,CC��ƍ� ӭ[7	�3#0�(��y��I�<�D��B>��V��@#֔������V�/W�t��p�KdR���n��u#F����?��4EO��?��$ax�C@3N�c��ϻ��s/�n�4��*y������y��2=�?�N:���8�(*�o�Ra�������1?U|�Y��`����@����>{镛ñ��pZs�FN8T�
WiN�����!����+�9rؙ�n_�c�C�n�僆l����iZ���{<B��	��������@����ˮ�~��U�?�����~fΜ���>5ʫz���
hwpy��`1���2��Ԏ�0a�w���MĞ}@#���|R{��C���r��x�@A�Ľ��,�@��f��?��=C!�B"}���L�z	\n�;5q�9���8;�c���1�L
�)�@�ғ���X9Gp?p���Ӛ�����lٲEZ3*++�Y��~����xhj��$>\���O���}��Ih`ί���uAhȻLv*�x�^�͘q׌/ڟ�����zh�'}lv:�9�����2��	���,���O{p��Ӧ��V��l�Z�����xp|is��l�(b�"(LQ����haD#�;��o�a݆]�&'}�Z��^j� ��;�88��E�x��\VxN��4k�|�&���q�[<z���&v�ŭ�*��_WVL�<c���83�N��d��蹜����o�z8Ys�!��̙3���z����w�}w���>}�P�56�W�rVL�3�#�[B�e���ZZ5M����� 4��@�y�`�'Vɺ�ţ]j巒d�PǬn� Hm��)��!���F?6@��I2���F�&xSS�O��g�	ؿ���g�(�!4�n�C4,� ��=� �����9��Os>9�\�����5��Y)Ԑ/`�/�]��+	��b+�r���L|��As�Oû-��<�vWuuu�%3ٍ�M�T�n�:���[������#�t���N[
���ht����O�nv�ޅC�3MSYt��ql�<��)���99QZY�Q�D��1�߾��{Ӂ���ҫW�` ߑ6t��}�?�� �Άj,Q@�,�CHe�RC�G��w}����A�ܰ�-���;��#^}��ǡ���T�t�����	 Es0Y>p��c/n!��n����}��W�������M��}@��%;�Y�\��(�p ,��]� ��RF�7�a ��L��n��Q^ؐ��"�e	*ds�p�M�Z��Q3�����Xr1�'�QK��M��|'8ӟnk{Y�N������/�$偉n�/��I�C�1h�4���Ǳ�?<�y�f���ܹ�w�#�����\���\��)Dii+�n� ��@y��P�8�v�9�N-9�o�{���[� ��z6��z�N����ߘ���~x����Q��2O���i�x�'�2䚂
5\1qrϚ�o���T��5MMC<�|B����Td���M�ܢ�S��Vz�����}�/v|��'gw�r��&��b
0ܳ9!��)�	]�H&�^yѽ�~מsϴVgDnݺ���c���Y3�0�b��ˋ��n��D���dt ����I7?ѧO+�e��?��������m��*�ez0?95h �e��h�9�d+7d�ˇ?< &0���c��Xn.�X�댲�â ��H���6�}�L�v`nf=��D0���䄑��4t��I��� ���.�Z[u
>v���t�� �ąLu;s� �a�͡q    IDAT�@@����C8���9�ҥ��{�3�a}��c�h��0���	^���T9�M�=O -+s��v�P����	��-?~|����=8x񫯾Z2��;'gt�"S�B$�����������c�`��B
�]3~�{�_��S&waq2�eu
[$<3ъJaD��7��J����z����Ҷ9��=m���[R�p�N����z&#]�t&'v6%D�������N�3��־wW�~���;g�K�ҿv:܊�d1k�brCI&ӹh4�Z߾}��v�m���s�;�Gn��/\xN]}���L�T*�@j]�$�LӢ�a�ش-��L���ɀ ѿM��B�@H��:��1��"�Y��	w<�����k�L���	�xg��>4�m�=g�t�������O��`�d�c�y�#�v����Q8�k�$�l�v�?9#�u3�-�$��8�k7�v�޽����c��X|���鞄9�@�; ��Z�'�	����A�I�-�u�ܟ��;^rɳh���;�R��.8���~�������g��X����D"~�-�|��Swuța=�:碲�����՟Մ/���\*\Z.�"�����v�t�ig<���]�?ʵ)��d�7�|rp���&Es��3���g'�2�h�gDM"-�A����7^6����b��Ν~�+���$�I��6�	�rֆ��l��p�����_~�����In/�������'ϊ˫��j���͇���@z�I\��]N	���-Ĭ�d$���: p 5 C�x���1�I;,�&͸h���!o m\۱cǖ8o�k$�I-3�����3�i.&��N��k�Ih0&���i<�?� p�l��H����O��/��@_�॰� {�N�$�3v��{�CY�	@G;�w���KK
���an�o���N;� �A;(G��G}��L�ߟ	���y|��#F�x����=̴7����+����RN�f�R9�sH��u`K��;'U�<x�����с�Npm�|gYJ?� g@���a���E���"Pj�X�Jc[��{��x��B_kS@����ek�|�p2=Г�wV��!��"R͚h��E�!�X��j�Ov�7���eÆ�I���YS;^ӵ��tEqZ�W4ǥ�������x㣏>�\�&h��t�W=|��G�]��Ԝn��d��֙^; ݾ�SSU+M��K�;@�9OE��;�S�#�@a�>f�:�B} \��ؠx�	�D �=D��8�w���ak�.`\�#C��&s�5y
t9��9�u��)DP ��$p4I��8h] ���u�mc(X`�.//�DC�7ڴ[��@;�㫯���d4�'ä5 4�x%������S�8)�H�d>���ף
 �>ě��{��5i���kv���^a�|����c�O4M��x<^a�	�o�# �m�液��[n�q�Å���3����[sK��"�p*NM�������+*fIT|��)�s���/�����M��y�z���E���׍d2&��0���!-��U��5��Ň����.o}M����)�(B��朖��`�'���~��N�鰉'��ʹ�}�<yb�Uo�5A׳��5�Jpf97g����c×�����X�Z�0�2 �S�f�:O�$C��`l�����&��͹���u;��!V<����i�R	H0�(���-�e�rf������ڨ��V�L��D7�8}��ߓ����O4���0��}���~k�<"7�;�\Ih��ly��bq-6qjXԱ�����E���/0�Q��XY�Q
(k�P�:���ev@G۸�3�:�ǳ����q��y�w�Y�1���/�/�h��x�`͡��A^�L;��+�w�)�́-�-�j��E�/��`��)T�!¾�t�"�
�-f�Co��v�����9j�k��M�t��0�7ڗ�ΎfE�/O��x��##�3�A7E����1=�/*m@<[�����\��#B�#Ȧv�,��������o�7^۩�������ŋwx��e�v���u����ʤ1�� ���ܮ��k+�׍��iM�z�^�8j�e�@ �͞�5��p !� ` ����eR�yS@�v��qIeh���4L)�0��ln�Oa��|O �c�v�fi���>��j���j�y ��v�-� @#�2�k�t�:C�0vM`��pQ@S��ߵkWi��p@�;ޙ�cC�8ԉ������B���w�����9Q�eK2����/^p�e����<���RĤ?���{�.��d� ��@��}�{�:�R�>�g'1bD��wu�[׬�4mޅ�m5�g3�BC����>)�K�e�Z�˱M�\6���~ZP~�6��7ߌ���#��;c��S�_uE��TD"�MiC�fQ������5��ծ.-�d2׌�j���L�hZY0 sl���q��\��;V^��SO<�c�j�N�իW�f͙������z�2��N����X��"I�SU9�vM�vK�n���Hŋ6|B�}�dW�x<��5�r�С�P`"'�������f�ɪ���7���j���n����	�v�3���e�Mpcx�3�ù��N���ߓ<G� >7��<P?@�. 3� �6��A�Ƶ� C�Θ�w�yGZ ���4�S K��-�������9�6���0�^
Q�$����������À�����k�&����W���,[��q�a�Xk�O���S��g߳��ܘˆ�<:��W�w�3G���"c�[�����\:W�&�7�ݫ��匟�yd��m�_<�P�/^_��C�8ÝH
��-�S�R�HgDSN5Z6���/�����%��z�lڴ�f��9@�4�̒�+��j���0L�����O�ِ�nk}����
����/;�믿�c{MM����eM�T@�
#gŬ���� �2֦M�3R�B3ǆ�?ħ3	
5Wj���66 ��A�)F1;$�1�A��@A�=M��'��EM�Y�HNcV9�C��n�Fg|�Hj�;5QƁ3�,u��" ��:)�ЅA;��	s(��!ܠ^���&`^v{�V��pŹf�v�a���h�G���>�Z;6z+�!���I�\,.�Ǹ�:07Ҝ���B$3������P(�뛝:u�yѢE-��㿫'�V��O�B��5
�5�}!��v$\�CW^~�-UUU�ʹ�3�Ɲwv���7(I�N-�4G��)�.Պ�(.�};�T($�U�g��>���L�6�US�������t��+�n�G�A�I&E<����۲��t���__1���3���k���?��|���+}�ހ�Nm�V#7j�����z6b�M�sN{,�\�9s����˯Lɤ3�������q[Yɐ% @'�`�f%�q�5�9���4ɪV|4�y(�@��o'�QS�`���Ʀ�8h��ΐ5�ڦ$K65IС6���)N���khu�{���l\K͓@�v�e�tFr慂����eB}yb�|'��D8�~7����"`�����5�  �|h� � �E�-���Yc�?��Y�(���,��c։m�&B���ܑ�Ǳ@8�p�L f����5c�q�7}�ĉ��-�~ٿ��9s����V��r��i
������/�5S䄞����Y�<�!�N���[�lY�=>9���\�lN#���'|%�"бR�E!���x/�s�k<���w���.�&���z/��P"���/�9��t[�Q��&�Қ���@�{_TV�p�0Q'�x}���~�{�4���δ��L�?ǆ�t������4u���z��i��o��������G������
�i�%���o C�  �F����/�A��k���hԒ	�D��bhs
�A�WN?<�f2�N���2�l�G�5���h��y��1&���h�9����fx�4��)�0,�N��o�e�����/�7� 6��SƸ�_;� G�q|2�>a��C@[�O�UT���C�-c�xH���/$HC��\ƨ�7�yD}���Bם� 
,��^h=!!k$��7.�{��A�j�O���κu�7�s]2���f���tw t�{7����}���w���{��j���\q��u���t�ki�a�u��7���**�P��%�I�O:�1��?���{U� z��g"�,���h"s���x� ,y,?��Ȉx&+ꄙl�z�/��ѿ���R3n��So�O��4����F�H�Ch��gu�>G�={���;��;�]y��>_��L�b���;�ҺU/�6�X��c���	��`@�&��%�0a�/�`d'u�����M %0X>��"�-�	NA��f��,��8��8�i��>�����Rk'h㳝�λ���O� ��#�k��b~p^X̏ufXj� k�'�!_;�0�c=�IA��o��~u��t(/���@Ȳ��M)���������:!T�����Աd��O�v��gh	�zS��Ѯyv~��p��u����_������v#v�ǭ���Ŧ=����3�g�9���G�5�Y���}و������D�
E8}ͭ�.��r��|����g��'=-xt������R� ��G���Ko̊��ߪiMx�n��(�ZFd�S"��E�C��;��_�9��Z{r^~yE�ܹ��WU��P��&�`�a#�ǥſ9>uw�UWLF�֞��Y��Ww^���.���L&�2F��,��-��~d)���2��d�cC`����,ӻ*Cq|��b������;�
��PǃX�%SC�AKd�9��0;��������E{���^|OS=�O��N��&�:x�����?��uC� �<1w����Wn�4�2���H�7Y�L��0A�3���d�k�0 �|ݺu'��Ծ+*;�X^�VF�]�VZU`�>�xB��>z���g��0��>�ħ��sa��|�����s-=��g��{ߝO�U���,��C���(.�]
�M��e�ٜ���7j��As$�˷�]��/������0]Q��ؠ_�;t��b�E�b���j��#:��_'��	���R}h���e�GyҺP�.a�V|q�)!���P��*Jo����?(g��i{���{=���*����2/b��d�wee�3n��Ň�Ie�?v�W�ʕ˂3f,�D���d2�/���B���b��Ĺ!S;'H�>a�n�$|��쀏2�4� Gl���ivƦ?/�/�20P+�_��k����:I�C�?��:-��H�#��v�/�J��1V�8?v�:Y�t9�oO:�ݨ���~YeX�r��x�,}c�(��`!d���~+��� ����[�*cN �A��YW'�#eyM=hq7�<�E�XC��ԉ��8�xG}x�n��r1��ay�nh����������3�<��y;���^�+W��̸��	��_nFk��Ϝ|��M"��	�4>>��c�w��2��<y�����Դk#�dǩF}���������[�Q|�ͭ7:W^u����)��ïVt�\��õ�]���Li]�YCx]n�s8E"����5fu���Z��c����z&'��'�s��O>��0��O�Jh��Ί#������ŋ�Mr?�>��K����ofk��7�wIr�b%�	�#�/ק�TM337[l�X�t%XC ��7�Ql��ХY7�77tl�d|0�9�y�-3����C�R�`F9�wӗM`�gf��H�2��I��i*&��B�=���{�<5\���k��1y�f� 1�
$�!)�H�C8����o�� 3�ǭ�yhjhh���)�Wg�t��s�(��q=�F_��ݠ���]2�v>E,�L���f���$r�(��=�F_���������c���k��\���V�m�i�P
�1ɍ�LR����y�)��\?����(��Z�_4藾-�s�������(����*Be�_�I�4E},�ܳ���+}���%��+WFV>���4�_�Kd��lN�ܪ�S�)	��Y=�]u-���F������ׇ�O�u̶��G	���掄&��c���̜��z�_�����6�?�?l�@摥ޘ�f/���/Q]ց%���{����A_�O Ч�����D3�=�@��c�m����g8� Z&�aQu�w�-�� v(�A�#��u�Ϙl�k?d���z�4|���%5y;@����\�̜�$R� ���v���;���3cC?��B�a�\���zX���6��a�*7��|�\�������I� �
s��)|�,��w��׽k7Y�$�� �(�8t��!l�G� s��h@�~�.�Ac���t�<�W��6���}?�IڻK�7��;o���4��PA��G�/&�2Zz�W�|�)�L$�S�{վ�΂
M?���!����D��Dx�K���<��������2��W���=V��+/�S���r4�]jN��#RzV��I�k��5sM�a���/�ݔ��Z�b�9s������YC�vN�ÝG���?:t�Л�9�v���Ia9������vZss����v���X�,]� 2Td��fgd�<�&eu�e�9�mؠ(�F)�Rl�L	
�B9��u�r`s��h�$�� >��	(�?�6, 9L� yZX>�}aB;��|������;1����1n��dg�6r�o;OD�p����A@g�[�b,0k3�.��Ü0V���m�EϞ=E��H.���Қ&�nݾM�1]' ufc4��J�f��-���/֞�HF'P�C�d,�G�ᅾ������R	뙢���#Ѣ�K�>����ۋ�3�lٲ�EޞN��(��2��v�%�Ȥ�N;��aW]5�`b��}���5�V�Q�ʜ]�уAʨK�,/�h�pEJ�6!V{�1�b�����������8xۻ�?R!�9�BU�2�);��)C�WEl�/��r��{���,]����K~����J#i�w�M Z65UU��q�7<p�	'X���.���Y�:=���;�Nǯb�X@�L��fNiP��w֐�̷�*�$�"��foՉM�36u��M�;�u$p�xN�A��Y�@J�89h���P��vI4C #�����0yIZ8i��3�C�Ԗ�6��$��Z�ۮ��GNs5�g"�G?h6��e�GX���B�m��r
��s��|�� 4�����I��++*d�vj�Y	�t���܈��N�BG�!��޼q��`�Gy� ���� ��(��s�u&q�i��<�9���E�ȃ���4��n(��.=l^h�ʕ�9��\���TmF�����{�s������#�t�͓&����C^|��hC�ZE)�Ew�n.��P�r�t[s���~���{����ˠ����7���Y��������{�¥ �SF�S�hHg�%��W�w��m"�t��#>���ǌ��Sq \ʊ�ŋ�=���E�=�Y�h�+�@v(�綥{k֬qO�t�y;v���x����h�@c��O
=��5~�gl� ��y(5d��Sج���E5Yh���:(��f�����:���~��g�JGw� ���h��S�i�~�gj���	� +fy#�ۅ�F`����|�	�	[�Z(8�����Xq=����O��~29��<��n��X�J;XIzjjd; �I�f����<�+��33�1,������k���kt
���m��9?�{���ɥ���e%eeu:�����(����ϼ��<o{C?�����֮]������DR�{��,��O�4����Ӎ�}������xW�qp4��(Η@~�␈v��h�h����a��~��)ʡ��Q�M�:�?u��!�چ[<��"���'�5��c���Og̝.eU�O����6�U_wݰ�|�͆{s�\�Ħli]vGU�U}��:c�oҴ    IDAT��:��������W�yo<;)��x�޶�eN��-�N "x�Ǧp�f�|h}�<`�|�dk�=&m���XP��W4)����`nF;����}���/j�/�Kk�@��j%˝��K� MZ0�����m��LfCB!5\��a{4�1�T0_;�ȴ��m2Y�5���6d�#�c-�k��1��x������ѣ���.���r�-ԏ��\�d�� l�I���R��\R��Q�@�����c��_����P�P���r�|�#'�w����Z�n�l�Ν��駟�?�͞�t:���h(9�w�K��G:��N_[Q]����߽{����0wr���-��( �e%"PZ)>��t?���cFE����ˠU}���G?�M�aޤ���N�P="�͉t,%��Q���F�����=c��m�cݺ�����k��Y�@�� �7o��|>����;��!CF�q��nz�Z����~�wۤ[.Kk��d�`Í�鴎��K��ЌK�8 �v|ƃ�M� �wfk# 39��S,@
:L����;��`�'{�Z6~g�S� �po <0&2u̤F �v��̉�-�3�⏠�> �h^���kYC)�''˝�u�!�@0�P��E�+���&g��ca\���),@��z`�0/~ � v��fy 0�`ލK�u`��rL��X���:7m�$�¬~$*�o��2$�a��g��	r�3AꇆA�A?�WZ�x�ʃ�$�Ͳ?��8�ǳ6\�q��k_���ʶ�C�?����?�5k֭�t����3�gH��<n�\ɴ�N��g�y�U�]6�B����~Y�;K��9��0�H"�!�<��\���p��"���ڣ��.���T[��lQe�ߝ]Ԝ��d���9�K�5]���39Q'���hx�W]<��g4��B�\����g�gF]�*�C�>}��;��4E"�%Ç_}�g�Y0��������5�w?��=�4OjhlvAc�� N@�b�-ֱ�����@0!� ��4+˃\.���ج�	X ;��@�r<�}B[ y��+
h� �n%S��#�A�@2�g���>�;��� 0��Z<��xy�K?Iq����� ���4�t
: ����O!��~z�1wp7@p8蠃�����PY���B�ԁ����q�D.C�t]��=h�ђ��#�:#0f�4����΅6��������$���ݻ���\�(P�!w��{�B��O�����;y�O��v?~��}�L�2e��L�_/s(g�}�����)��Ϙ��,��ʜ�����tڴ��G�{����Sg]QV]��T�(�y�������t�"rᰨ������G�<��mq�����Z�Wϙ�S����d?�f���.� -K��@77�TV5�����%K�t{r٣�:�1��/|9!a�V��Z���Ν+g�rˤ�{���~��.�J��'N����5!�uB.|�iF��W̆Fm�v-0�2�q�ǃ���0�Ӿ!3a~c�
\K4ʣ�7�|#7i�3-M���:�q� $A��#��!] s�����L/�'���<���6ƈ�}�<��+�r���J'У}2�i���o��+N�6N&�����mh��x���Ac�VL�
c���BƁ�a���Z�q-�$���M�d��.��#�s�~`��Og�_8�%�c|�`m!��=��O[���FL�ky�-y	�XPX¸%�_ϴ�á|���Z��?z�G��TW�p���?f��k�=t�ڵ��y�⾐�͠�%b.��-.�4aB��nݺY�"����#�_o��4�>$�N�2�*�.Sz�c�p����Ǜ�u9������P��q��
�/�~[׺�͉�Ԭ.� ��"�ʈL<#82��}<�K�[0���X�3���7�P������I�|�����o<��,x���k�2q�=�\��^�0�%�I [�:�s�'��G^�S[���Rd?M��R<#Z6t���C\��� �; �b�F  m4s���3� P��(������? ڥ��@̳��Qu��U^�/�A�&Quп��5d��ba�
�r(CS2-���+�X1
Q$�z2�If�w�u��a�1�8�e� �̇��>/$�I�y(l%�1�CX$(���ˉ�7�n�u�&qF1�}��a��ºa�%�д�L�����>6Ś��ꁵ�!;�p�TH����t����b@è�F���{�awL�0�fמ��R�n��bŊ��\��<���Xa%�U�4ͤ��Yt��1���ӧ`,�/�vg�ͯ�5�$��eQ<�,����eO�+BE}A�](/D?���9��rO��
��U�;�hC͜`s��[�6���!bIMdbI�)b�"V�{�1�Ok#Bܘ1�����O�;JI:��@�$h%�V���)^�x�1�M�<�`R�dW�}���.�?4�H�����h�,���i�ͱ�Z��?��0�f�Q-35� ��;M��� ��٣>^�r� 0  0��ϸn�=�
��u<�������>Cc���F�>� A�( a�	i����� !\��Y�b^S��������,�e�Զ�!q�/�:C�8F��y��y�arG���g�m2<�Ř�L�`�اs9�-$N���l�l�*M�XG�7Ǎ���\�Ƙ�hQDjബ��� � �>y� �n(�ւfw����������Fd�Y����=��;��'�\�+�@{�?y?�-��]����`�.�Z^2�p8����0`@��u�h��ѷZ4.K.J$�;��?��N��|���3�+��"M0"���X"�$�Ċ
�*QT@l��ET@��hlX�Q�meپ�����s�Y'�}SP1q��g��{�=���y�k����!��r)�� N_�ԋ�E��tZבC^2�A�����9����^���s
�ڮ�"�JB� zk(,����o�8_=`䰋���{��۷�gϜq��-[���6W8���R%-"t���^���ѣG���+�l��A��+0}���{�����؈P(d�t� ô�� �ӻ=�It����# ؐ�!���%RJp �,�I�2�B�CY,J��~�����PD�b\O��r ���;��!-2y�ۜ��;���l��~ ��@N;2̋�7����Ep���%uڇ�]���=U�L?�,o�3�߳�1WJ�X;8�A����1_�m���t�������I��Jj[�oS}s�1��� 	�|̇1�^�f�H��0�|{���|0G�'�88w5z����3�,T��L��9��ð<t��w�������O�W��X�d�m֬Y�E"�c�X�b�mv�|Ym:#$�^2���a����+'�7�-�g������O-h�(�Dz�Z��U)�U�/E�ś_"-bi����s�	s�޽���w9tx�o~�����.t�E�=C<n��̈́� ��5!��t����3N��G���C�}�ڢkg�|c �(���sH�x��P&��6���/���3�8c���^<�>x�9��u�%�-5k�f68ڎ�����i?�78����:���b*L�k@��m� Ȑ� �!ޜ�P���.�F�+���IK�� 1��� J� �Բ����saX��謇�SO�c�OI�@�u��6e�#�S��_Fu�nw�\_��,�B�	�p%]H���h�|���������������;7�N��������X�͛7�W��f�0���}��h�;�8�������p���獪x�^P;�uP!{6#�v��V^Qz�#�<���n/�.���U���k1�^�3��,OD%���ݻ�E3g���a����^6 ����*"��)q��
��%~�Jie'I8=��h�ٮGu�1j�w�9�M��oy��Y����ma�K��[$��K+�=�S�bښ��9�ܟ����[���],[����w�~W(G��ӪT��N��q����ĉ'�p�	?x���My��;;>����ۂGG�Q'$pm7���9	$:6X�TA����9�Y�x���Sb�Z ��!������@�?�(}S*8���u�O�:��"�	  �!f�u�0C��<ہ!c�&�P)���:q�g�A��ȶ�SmO59A}㾩�g�70T�sJ���cޜ?Ӻr�逆~a���X09�C�P�cn�SϘp�3���)�L��ĵ�|���[1���Y�0>�� �=�����@8 |�%�s��o���L{L�����X�o�v@�8�#��+�4o<�W'?1nܥ?8�~K=mڴ.���#i3=I��/(�8@&C�6���3'^u��=z��y��zKo�tg��w�L/jl9�8���̴��]���[�/��%�tKm,��dȀ��N^����7���/{�����}�HQH��#@���$c
�����U[Y���;���A�r^�p��k}x���D�8���*��.
A�߿��믿vȐ!?8����v�g�dӦ�����$�t�=YU��L8>�APA4A�A��5*@��c�+�35ոhbL�1ydx���� ,h����E`�o������G?"�>���,��	P���3���N����amx-���?�)��h��FP�o�V�D����i��g��e���,Q�N� �hO-���!���qr��H���%c��ŏ� c�aO����g�|�V c���A���9EH�8x`{�Z���-����^�l���tVg�Y��ɀ�#��j�F̴�j��}���{��M�������Ǌ'��x<q��jubO�tA%�ς�֘�n}t��	�۟�o�K/y^~艳�_��P���)�ynqx��/��$�͓��Ygv�8���cZ�؇�������\�~�?hv�c� �ؐp:.�`HB��4��M�NՓϙ���ahJ���<�m񢗟L��Ch+�ʝ�:_�4�***����o�ԩ�w��/�K�W�~�gJ{�Y�P�6��INoZ�s��HH ���㨣���fr�����L�RU�h�xrڝ!�A�J���q&  � ��L�?^�4^�1�J�s ��?�q��_T�2�%d:�a�`4l�0��ɰ0̊.�1[�ύ�� k�ybVZ�;ʠ �`��F���{�<�C;6fR���� [0XP�Ӧ���o�?��0k���g� �ǵ`8:HE2)P&�#<�ͼ�٪w�!����_*F�a^|0�Kg�ZF4�랙��r'�E@G?P��UPP��b�O������1cb{����dѢEEsf��]8:��t�c �c���f���d��=Ҙ1cv�OK���Ko�voy2�Ǘ���a��*��)��[~��Y�&�����%�;s�Kn��_j�����} �nC�t�}ƥ!%�Y{���缽/6���h�GL��G@G:�.	��b�ٻw��M�6���&�/��}cҤI�\��C�@p���̄5i9S�R�I;�ۭ�^�xB����/�V!N	���, jH�5*�I���I��^�@�_�g{�J�H�xG�EY @LC� s�dp��P�s���/=�� � \�'^�xN蟒0� �0���<�Tǳړ�ҧ��� m�d��xg�@4��+�f�[6����3��ǋ���q/���F q�9 �PǣO����s�����ע�8@��!0C�Bi~٩{q���?0����?���A&�P	i-�J�?���aw��1o��fL�!�"U�ׯwN���	��M�nw�J4����L��Ŕ��f���?}�9�\��[��?7qrצ�V�[����Rv���C�[����rq��I��Z���x�A�F���N�9�7�O=�R����-����ӄ�)�T\јD�)iH[�9�Wco���^^����k����M7=�J��P����� 1���C���[ny���+(�2s��5�4N�UV�=㐥� �J�VP�މ����K/�T��~EP��vP�A�K+<���i�կ�YzL���� ��! c�k��@�����Z��j]\����R+����|Gm�ࡗ9��wclw6��3�`r���xj������� d`* �̔Go{����������X��e˖)u7���`�poXW�>`l�>ǽ ���ˡEc��b�eOQ�}0��wjzȴa�k׮Us`{�6QL�i0& t�"���3��iMf�A;�>�}��p���}PRPt�����辠��j�3ƍ;u󖭷��.�q�����Q`��vۗ�����ۯ��ùs�W�}zFA tzq4]Xd���f�'�-���T����L�2���'u���p�˹�9{�r苦M:�]x�����&�n��"Ii�G�GSVi����r���������@M��Sv��}o2�(�S�M��e�m���ى'�x֤I���ô/�gO�x�G��~z�ݱxtt:�v�SZeYT�n�C˔� ��P������S@3�|�N�s�a_ ��W�=������BN���㻔@�5k��=��+�,p�6��R��a��4����6�Ƌ�h/g�6���cz�y�<0���`��ҧ��H��2�����,ǽ�V��;���H�C�p�s��aE������c�!ELq~Úa�X���C�:��L�B���q����kO��v�[0u�#��9���%���583�#V0����.��XS%��=�Ta�c������z7n�Ϟ7n��q{B(����/�����W<�N&T�ȓ��b^�Gg���*��.��������_ݚ�~���\{���隢@�[�a��En���oE��f[��{�������W����+'�n.Yb[��Kc��ᇍ�P�'���P��p��F�K��-v�=O9Ⴁ��s��4-]𫋚[�f$��B���U	������?��^x��h���\p�G�[����P[��t&��ٞ@��e���x<�X�#G�ƍ��;�-�+y�%h��D�G?���?��C&�B�'�<�6����Ǟ3�
 @�=�@	��/��@������=��}QuI�*v:�Q�e�5�qņS*D?��1_TSS2����Nxt�#@{=�i&�� ���u�}ӻ��A �<� N2�� 0�$�|� l�#� a���3��~�o��:�[9�R��@�:����!�f��u��)�=��^�,ڂ��S��J-���4�Df
s�� FR$�ɠϟ�l�~�����ۑ+Tc|�w��B#�n�O�myy����ym���3.�����J���=��[��=��uXQ2-�N��6����W^&�U�l��vI�p��G\�>t��o�b{�:'�^��Ǟ5�.8����h
8)q[-�H�$����T���ze�ٿ?��q9CR�7\7���ib,�1��YH�� |0a_�3f����ٶ���?��3c��[[[��%J]k�*^H*��S�"ܔ�@4� �����CU�g8<Д�)偘B���� � � (H�`�������!�1�U�T�*���o� cf�a!��5��Zq��2��� K�K�j�;m�x's@@�$N���� N@���-ݓ!��N�������r @q�\0ZXg�I-�T���i�k�B�1`�8ĕә}`�=�p- �ad�^��{�~�Ʀ����:���>�; ��/��9��0G2\���ұ7L8��(	���{S��&����e��>...�l޼y��������g��p��3����t:mV�S�+$t�2�2,��.�쪙�z�w�����+�fU��[7VG��h�Y`�ćT���RPY!���ҖN�3��``�K;�~��}��9���_�_���3���[��p^6�b!i�'�%���8�~�yWp�Ojs}�+W�,��[o����q�R�ھ����YXX��W\q�����ֵ��z|��}�њ'����d256������T���ũ=�)X��V{��x≊�.]�TIL�V�� � �tP�Ə�    IDAT�T@p�����O�TG�Ę�� 	�8
��҄� Y�� 1���g<���e��16 �R>�О�20�`azW�VM���aJ�١pٶu2�l�9��f𙚌l- ��+������@�I��hO5<�!��o *��i�������<P������A�ƞ#-/2- {�%�yÞaoi~�>��P^�Fcb�c:a�W�i�hj ����5�;7f��:��5g�'=|���<gƷy>��.,��]�����~n�X<��S�u�����MIͻ��_M=���U���<S��cO]V�_��PQB��!�|��K^Y��A���xi�5]O9�)c:W�з���hݳ�\�J\g6�]�dZ��^N���KHSBB�n���O���Σs�i��n�=���d*}Z,s�aƃ	����p8Q^^��5�\s�СCsn؟�5����0tŊ�����<���%36]]Y%iY>���k�?���w�QD�@C�2|Gw���g�}饗�@G&2����wc�}Ԍ�&8`�J��5 1��	����%N�r:��0�l�0�v���JN�~���k~G)�6ٿ���g�T��! pg��ﲁ�0�t�' nԒ�X
S�b=��F�kLos���&k�~�	��И���u�8���f�$����!)C��f� ��½a�aC?�k@��<��:�!�5F�W���Ai`���l|Xk���X-���{�U3g���������?Ο:e�X8|Q2���d�ߟ��H�i��tr�?���SN�̳k���_�غ�E�H��tR�S���+�G�O��e�*,�lM��{�	����˵��r��^z�d��&G�W�Z�vG��Ezk$ -q ���=�ҩ]F�ص�3��K����w�w��j�q$Q�S P������x���j��ɓ/<x�w��ook�_�2��f�ry(�*����^m��&d�q����D�-�% Ep 
�=^�hQ{�Q:Bl@d6E	��^ M�66@/ڡƬA����0�����? ���A�d|pf�6:�Q� 	��p��|�=���~ �tZ˖ʹ��^�ْt�DO��F6�Ai ~@��� N"[�G�y2�'�����u��a=��aO�.t`����Æ�uŽ#�k��&�^���?�O'E0`� �pp���:���A[�F\����S���I3�c��ڶ6�������@��=� }�N���wق����ɀk׮uL��o.��]�H$J��}5��>`�u�f��Q����BװOM��s�;��J�GǢ���V�; ���Zee����բA_Q����ӷb�sqNV=�|Y��oM+'ǧ�" �k��d ��Xi_[���'����U�sf�U�?��6�}t �����$���Y�����Y8eʔ�0`�Jj��}�&}��������O�w�ͮ��p��еT{J�3Q�(-r���+»|�ru�g��8S:�)����7N^{�5El�m�HGF�1��Z���9�k����&��Y����|fc�r\� @�(�1i�DNPf�9�i��	�T1�Y,����l�v�%;��d�����jx\�y�kk�� ���x� �~ b?(�cNx����1>�`��`�p���!��Y�u dz�ӹ{���X�����X@K�=@[�ϱ����}�@"Q[�=��/�aY�pP���p8{�S��Y1��d`�G��b��ř�<��7��͸SǝT�{���t�Xl�,����Xw�L�-�4��˯�j�7)7-?x��|���d����C�)S|^�xˊăҿ%�R�Hn�UV��>��o�+o�� ��g��-]zK~(vN�5,��CBo�*	���h�><������@����=bw8�mmm����6Ev���0�`�Ν��2e�o���_�nrs4���k����e�>�3����6CrR����	^ \�r9d	*��V����AtA�AX	6��>��ce�ܹJRă"��$��+��"�_H ������q :̲�>��o�	Yh�=�B�-���&��`�Egl�� O�@��gK�ـ�ue_X?f����B�$K�;��mtD���_�#C�`�^љ`��+L���ڂ1�B�MPS�=(3
���{`xU�����+�����|0iA�5�q�𙬇����%��u�B��E�RD�����Y۰�f���O�81��!����~�8��ظ�˹�at5�ڏ��u�ZZ�2�훻��q�u�ݸ�iCPI��:�Z�krq��c��"�����Oi�x�J�VT,a�7��渻ϩc�Y��� ���"t��%|Z�5���f8��܍���{N�rŝ���<Z��s~��p�q���Ū� �q��{��OΜ9�w���9����x��������S�N�s���E����fj�8$t:��)`��H�;t��#F�O<ўw� �/&B!���B�;����^�Z�Ş<��t�:J��%$H��� ���}��N��R"%t��� Q�/�:d��9�l�t��~g��W��z�4Ool�֡_~�:�����j�.���>{����z�I������&�b���^�x�B��p��{����A-���8Q���g�4�z�e�'# �Ö�yb|�qΘ��$�#0�:�>��g=s�[D�������p΢�����aw|��n�u�}��o���2�+�����˖ͷZ�}!�㬕�+&:Ή���UV^1����S�喝��Z�?�v������;+�#�	)3l�Y�V�E�؋��,,����fр������u�b�s�?3�c�O�v�O�7ŖJ��f�D"�$��dRڜ��hy��O�b��u�I�s�z��;-~��ǝ.�Q���İؔPG�^�z�7cƌ�kjj�iB�����z�ڵy����_~�e�y�7M��T�E�۫)2��E'-�t�;���jU��q&@�A��%��*d|�=��3��W_U����)MU7�REOU7��.�r͚5
�1&�"��T�c�t�ø��I�E_ L���2�h�(J�ٛ�$]�&�U'z�Z�^�s�k����̖6$-) YlV���MS͍k�:��vw̃vh�%��k���d�w���8��q���?�c�����\�_XbLSϞ=�T��1�r�g3hK;:59��ǞBs�1��}a�|1??ց�m���� �)��=.m"h�s��#��B?���n������nz�G�?�v��eڴiݖ��֓V�u�b��P�����y�������}������w�K���U��go�N�������t��"�v[��S�UJ:?�J��JJ/�~�}����&9����9�r�����񉖰X��n��@2on���"��mw�����S'�W����{�]__��<��5���M�~]��jS}&�w�A�����������t���l�v�ڢm۶�jk�w�����ݻ{��ѳz��������=��Dı-P���iL7ռE\s�e���?��ڰ� S��w���6��pH&���+B ���7�'�m�EI�Tc��a�
��
E�*` 3� (W���B\��DEs�� Ξ1�z�m�U��?�{]^IIJlv0=��{q\L�n�Uۅ�Ju?!+�_Z�fR��#��!��x,���*f"Ӟ�xb	�+;��*M�%��.mj���hW�����@}�б�j�T{��_����A�U��"<�q&�w�vH�5aZ_Vn��9��`ڰNac�����iK�����޽���j��q~�c�;�5#ʄ��@��Z㢝�'�N��j}��3O�y�)g�W1����g�x���s��}�0���La�K�t�BT��L��͛�w�}������>�/�qۯ:4�)GʊRi�lb��+-���*�x�%bq�"޼��G�����r�9����ں��{=��Q�ֈ���p�%XZ�e�,�]��n=��J8 ������}�m=�^��<��9H�J93^�6�"xxè;���gL�r�+���w{zO{�z$ݩ��+زeK��_~�s��M#[Z[��R�Ҳ��B���+++�lذ�u7$�rfj�;�1	P�b.���w�F�RR6^Xs\i��"�����B{u;$=��0��g�	4U� ����+�-	�4�c���R�0P��	
�R��v%!2a
� s2$jA.{-g���
������<�cɘ�ע-��p8�B#Am�P�s@�\��{b���phg.0 ���׀k����14D��xT���bZ,�M�I  �q������ �ZVQ����� �55n%�c�X?��u`��/���h��� �%��1�;����6m�7��E_�� |��?�53�qy�P��ՠ���=��ڙ�ݖ��l�yՄ	��g��䱘;w�=�Tj,2x�U2�T\��i�=�{/;��Y�j����ˮf~��=��hߢX\
]Vq������[Z"���7�qz^-<����cs
�@���ǺE�r��5r,$t;�v�[R���K eJ��^kv��=�K)�*��ϙ����ޟo�� �ͭk:�SJr�X�֝�v�ٳg?m�m��ݻw��ر��аӻv�ښ[nni��D:Z,�NV��4�J�(M��4�L���j��#i�/ $���1�R6��p@� �*-eT�O����ǎ���h�!f�2�?U�T�������e;�iF@�����}�1 � z�c�� �g��ف�*s m;�[abJ3�AB�R�vڴd�E���P�|�羡n�C1�Z#@	)J5�#UiJ,��UN{m��_��R�ص��S"�7�ͦ=�ʹ�]�^��;���o@��bHt6Tu�̇{�B�M=O����g	c�\@�w�:
���`�0.�?�� �`�xfx� ���۰7t��^����~q�d��=������ �t���w�jx̍&��9����y��;��ݺ��dΜ9?�ѿ��A����3��d��k]Z\�k2����t�"n���3�<����s��nC^����_z����Q��#�HKA�S�!�,̗�N�%��I���"PZrn�_���,�9��O<�=����|m�c��q�E��$�1i��-�TZ��ZK�γ��tѣ��o���W��d^*��g1�cO Tơi�a�~��ٷ�>��}�4M�ƍ�7l��߲as�ί�:����_"�����e�d��b����ժ@A�!���82��r,�s����$e�g6A�B� a��X돇�m��}A0f�y���4B��@�ѧ��@U3������̚5��"��jg����l���E����ݍ�p�CL}~�O���i?�*{�C��;�tT�1 b�����<��J[K����I<�ԍ�m*����w(<��%$m�"N�DR�<DW`�uZ���z��˗P4"�`X�E'S�Y%�|<%���X�1��f2<�ة 3 ��c��+f�搖�x ��ad V�*փ�w��16�$����=z�s��<���|�U���w��W0�0�����8�K:G�� ��h�N]=0+����9�].����~e_�#}��_�,Z��r���s���O-�k�; �>�,��ָ��z�gg�y�QG�_F}�����?��o�ZC甇cEfZ�\����.._U���Bi�;6;�~��/�zOr��k�����n��8%��+	��n��y�1.�� ��n�>p�΋�S}�
M� Й��j�n;�ï���Q�GgJ���6nܘ___�[�zyɮ�]�v�~ud$��p�j\.g�i���d�F��D�� � �+V( ����֣1]�%�t1�)��
��-T��6�m���Ơ�ׂ���;$<�	��V���� D��5 �r�i��q�N�m�0�}�X� ������~����/(����W؇U�2�U�r��ڝ�p/V�C��۩�͑����k���z�&�ծ��ذK�V���\ fb�bW�r:y�2g8���M @Q1D)����R�G#	�|dU�x"���]���ᐝدh\�~�Xm���q0�nf�iD�W��O�{V�����O���Zm��;۳�1��f��/��3ƂH�{���za�p?�EV�N� P��83�'3����a� t�h�rǞb>`J0>���9t��HP�T�+���t�%�=>f̘�Y_�oJ/^\6{��Y�P�gV�Յ�-*(ԥ���%�p:���O6����yj�or/0<r�����}ykY(ֻʰ�7���.�|��W�Iv;���ylu���8{�&'���Ǻ��\s��5vl��M�ɔ�?�d��kH�6�W�.�gw�%�@��Z�zՓ�x�����]8���a7�6t�W�|��H��B~��n޼�U_��`ݺy[�l�\_�02����Ý�6k��n/D�d�5���,;ԉ��\�{���HR�C650�xSu�V�Xdμca/ �xAR���̦s��ѣ�wz&W�`
)�	&�p/�~G�(ъ���j�V��	=����#��O=����f�1���jwn��f*v�3Tݐ��/�E{M�g1I�R*液�R�}����a��i�Ӫl�$ă��>�����L�/��n'ӓ����V����'�@1�H(�E�*����L����Y\N�f�º�xv̼��́��T���3e��{��q��{	5Tb��v��aW0N����@@����z鰥R�����pd���D1�}@z'���g�"�������>h��6�c�q�,�B����� x<��X,���~v�mg�uVΓb}״eo���O�>}F[[�٨���R�_��Yt��fI8�?�~�)�9��r^�����gw���_W����*ȃ��f��+��"qT�K��b�t�9�f����8�i�� :��c�����>>Q�&�r0B�m�1�%��z�Rg��xǏ/�t_�>���=���+W���N}���p�O&�C�6b��{yt�4�˗//\�n�wǎͥ[6m=���� �����ru�Z���t��DT���HQ-�p����& )~�:��/�D�B��H�
U��))ѻ�jTHY K���F5��i�$3�4˄1 ��?��#5��b|1��u��#��1��Ç�'��8�0@1g<�2��$��}�!�ꘪY��
�֙��L{��)MǢpЯ����w��#�XT�|�bXRbX���ҒB��,��#i3�|O���u���p�-8�5�#�t��HJ0���finH$�Pɓ��x�
���T}��ܪ�tG&<0�gRnj�A��V�b�jm
l�w�� Cu�0mp}���;���:���)x���@�ά�������{d�ڲ���k�LC���@J�-���{�zq�h�̆���������Sv��ӦL���?%�?\�W �ܧO�~Ckk���tڋ5%�C���n����s?>�ƌ��f�\������z��ֺ�rp����=q�y�SZ$��r��꺶r������7�����,XP\�ꮼ�������<������f�QS}�IW]�O��1�����<k��Z���@E�5XY��y�7�x���#��b����;vl*ؾ�vPccӡ���]�K��n�p:��v�ݥ���ں]�i��R v E�FqU�$t�U�}��8D�R5�3�@; 1���Ꮆ�L1ǃ
p�e�V���X<�\������/�K{;��Y�K���r
 %�j[�1��|�M�V'�V���յ`0�+�GF�װ�Cݾj�*57�Z�aÆ�v�=�X{.z�00�7�;�DBj�`�U4Pɸ���ۙ,eN�[D�N���)*ΓҒ|))͗�BDah;�ϣk�pQPjvC��W	oa	E`�IcҤ~%�v7IKkP"��ڢ����嗲�*I�Mٱ�V
��$�Hi�8��.`�;�	���Rs�)��%C�0_�m�� �7J��N+����r�q-�Ěa�8.����Dz�c��Щ�0Ϗ    IDAT���;���R:����N��;}1`Ơ��AIk��6����]8N�춥�{��>��;��5��o���/��M�4�����M��ú��5cf�&$�͒r:/�p☉�F��_��X���W��պi�	�x��|_������")��eu�Æ�fTW���	��X��*���
B�_&v��Dcbw�E,��Z�1���%^R����R5"�a	JB_��<���j<�C�mj ��^��C9�3g пs:
lݺ5�ƍy�7��ZWWwL8�eF��Ym�X�E�c�X�'!��A�@��C���()��!�J�+���y�q�О![TES��o��:�gw�"�^�v��W��P�A�S����:��A�� �z�l�;Ɔ�pE�T�*��Nm �SE�$6��qO8�UR����˚ ��lF����#G��GyD���v�,����N���s�4��H���0��� \,��R^Q&/��XEۈ�.��-ҥs�ح"e�ҡ�T�򤺦B���=ǸN@nMK�d�`�C
Da'��� �_���-;e�����@$!�PR

����I���%RT\��U��6��+>�ë́��sqI��t��:�H}_\�w���� �B�bF7z���)�� ������@K���(S����z�Y��2Y��;���s��4�1�f�c~~��0Gj�,�6�/oS�XTT��f���5(��U�Vy�O�>����R8��UA%�.�t�ӆ/7z�e'��:׫�W���Y�f���lٶ���}��(��Q
���Jzt������^ۜ �����?\yCa ~Azw�����	��4��HAἣ��xz�}P��֛���Oz��� 6���"��"��x<�>t��ٷ�)�;�r����.}����7�J��J�S�mv{'��Q�6�J)g6�Hѻ[����@����=qm�ZU�����鲕 Z��N�4։�d�+��)���m|G�&:6aTeB����ԵL�	BO�:J�<��/UH[�34	cR£��u��Sm��F[uh�7 �B>:�A�M�]wݥ��g�C�~�T�䣇j��E<J���$�����8_��O������(~������0���/�{u�����P&����s)	���UڸWV�LI�4�t{��42¥Rb�$MH�aii���d�m�y�.��m��[k%JHaA��T�S�X����$���D*�رJb��VG�
���,S�45�hX�>���5�0_8; ^�/�E��u���А�Ø���!CY|��
�X{�~�9�{K�!�8;�c�+�U������#��: ��`4F�y�f� �p8֝|�I�t��m^_�Ƒ#��<|��u��v/�@�'�#���_>u׮]��qF�X���q��i����cG���W��k_�㢗_����^�=��͗'�����b�u�ás�?_���eS�K-��V	E��u��fH[�U�CaiFtT~�ӣ.�8��1C���@|�k���~���I�'o :��U��բ<$6�˵cРC����[��&�|�6 �%KwZ���1�!�<yy&≢t:�귃Hf{q��aL?$H*8�70~��M�Ĕ@��k�D/�}bL��SPE�l\O9���1�$G��!<��>kϓN�>����I�?�)U�@�q� ��̊bX2���Z]gS��@[�#G��s��!�ԡ�@��#�ҥK���c ��S��Ե��z�x<y�֊�0:h`�p������� ���Ï���xEjwn��|�z�RTT �J�G�J�ޭFj:VIQ�_�|nmS7D���mZ��<�+�/ߩl5��4�-ZrO�u,v<��t�*�-�����g����6��M;$�0%��L�S��ܥ�ݘ�$�)��̓b�2��Je<�;Tf�cim5D�oOsޕ�`m�^hj�A�8����`R�,���-����a�poxWq���p���r)�:�*���)`q��S]ա��B�
}KtZ`���g�Z���N>����5V[[[
�6z�<K:h�ۇv`C����k߆�|Wm��{��W_�s��+�K�8����2t谋�����nݐ��ɇ�ڝ�7y��G9lN�t��uM<a����S��	�����mo������D�muH8"./RYZ$HC0,��t���v�EO�26�������>\�Lq�RICs�îly��G���M�2�7�TUUi/�}��
��7_�������r� 6C�h��i�Β���DR�ʌ&ډ��aL3�ր�F������E�9�)$%��C_tDRNZ5-�F;�Zc�M��b( �`��=.� �B0�\��A�dF���Ĝ�>�:�'<��K/���r�#~�^�1��H�o�92����q0_�$��|���?�A����(�u�=r��gɧ���d2�l���ҷO/�ݱI�}��t�P*>�S
�^�ڹF�k*�[�J)-����a��f���v�jw"}��`��o�����w=�/ |*%��# �a��EL�4Էʆ��d�gd͚���u���)(�z��M�wjOnh;Pf6�Rሸ?$��vF9UJZ�]e��I���2n��=����|�8?�jO�k��8aFC��c��aX����p�c�"������q�+`�1_���|]�'[�C
��� �2�Q3�)2d����x<�D(j�Fc��O+*+�r�aG��ٳg�� �> U{e �5�\sͶm�&�H~6��o�9-�b�Z=�O=�9ϰ�Wn,��yO�;�����5���*Ag:w������t:���ce��@��xI�g��qIa 6Yj[�f $N乵���1��X:���{a�E]}�Org���w�|��w��Z�([�iS ��Y tH�v�}W�~�n�>�������IA�7�x��՗_>r��Mg���$��2�V1|�6jJ$ .ڹO'!���%��3���i���C�O'$��%A�wt���	�ꐰ@�� }r>d�b�ؘ?É�	혟s�5��c�f\ i�V�6�U�l��;a&��<���f�r�g�&s�:�F�D�`$p6hh���2y�de�W�ө�B�8�ty}�*�B"�ŔҒY��B�)-�Iq�Oj:UH�^ݥ��Tj:V��m����SQesw�]��K>�#jנ.Q�\�J0O*�����LI*��㴪�&f�R�oڰ]>��Y��SY��1������.�X�v%�GQ$&��U�����p:���������^2�.ڐabdB|�(�e�_�Qh�NmN`x$�+ɘa͡%R�*�R���#����Sނ!��
�{h�s��s��������|��z��Uu�P���B�P��jm�z��[-��;V�9h�a���`����T�&M��u��	�a(	=���a��`�0g��#�������h��?/���C�ک�7��n��������[V�W���7�/Ʀ�W��ts�����ʫ�9��h*����y��Ο�k\��}�ޮo���I��u:��� ���+�Y�{��=g�̛(**�y�_|���g�:�b��f�f�X,f��9�hO�4��$�|��%2m����G�c��nTLA8�����	��I�+fa���)��lJ�َs �T��O�6֝�̘/֜D}��q���D?��T�2�,�4�y�=->����/�/�9����d�������#�{G��n�A���(c��G=�kj���|��R,�`���ԉÚ��]��{�ҵK��:����yRQS�$k��!�d,����)�\l�<pb c[�22�X>d��7�	|�I*�Ik�}ô���I���榀�^�V���L>Y�Y����tO�X�S� Tâ��)�{J�W^�N�Z�H(�"`��0��w e^O�߳���]�D�˪ҟkN0�Ɔ�r�7Cq�.�}��NOt��`n��Ff �N�S2�5Yٚ!�W2�LՋ�ɴ���L溪�
�P]�|P06�u�ΉQ�M<�L��R���XSݱfq�~�u�޽�o߾���W^y��;vL�Z�~�5 ]9Ef �鴛�tj�1ǌ����uuu����n׿���4ҩc�iN���0B��� z���k_x���L���O����
��LzS8�lrz^=��_�tv�P��ז�5��N(���r*[|�4��u���-��<���:����{���O=1�������XC0���ӹ�޻��:Z��� �:ƜjcH` ��H�"�~�Y16Im��g/U�X#�p��Ts#|�Hu'5 ��h�\@�!��������z�:7�O��� R̍v|\��!
 �{Vj�L���q�6�¼׭��]�Nqh�>���uL��-4�:�������0k��C�m@�/O���u�(k?])�����mҿO7�ԩ\���"]�TI׮�Ĵ����K�@̵�*�����H�b��u�S� ��ڟ$��쭖�X���T�tB�(���3�<�(�j�m��ɇ�T�|c���%%K}C��=~I��V�)��ՙ�hy�ʑ2Ov�ܮ�k�����eG<p��	�C�SPZ�y2qM4<�tl�>"�;�����d"�t�#H��2t�g��u t́s����S���m��E�n�ܥ#�/���y�̃���(�YXX1�!
oJ��'ee%ov����>�᠃j����������?~�]�����h�ϯM�v1�r9�t:��ȣ�_�}td�{f޼s���匁T��K�N�;=����dD9ts�v��?�;9?�+�}wI��M�����Z�!i	ĥ��~��O��h��n���CA�ŋ��P"?��-��PU�x�@=�L&ۺt����7�tm׮]s���k�U=���K��ٱh�0��� <t��_%-8t-g�:5�kչV��x^����Qr3��� b��HBK�7�)٢/HFT��0B)���bȑv�/�K"�51G?�3~Q-�>Ƽ_�	�
`���6�օ1GN	�Ap����}�vh�Ù��0,�L�� �>T��;��U����3v�E�*$�A?�/U�E��ӏ��-�s�ҳ[�t�Z%�zwW�i>�[��4���T��q@tህ
kN���m\E�������C0��Һ��)�z:����ZI��p0$m�qy�O���K[0$�w���CF=j��"	il�N�6�]�B�lj�ׯ_��{FC�Ȝ�ak�s		{
���S0Bh��U:݌O%v�X`���g
g}b�A����ؘ3���!��N����R:�{fW�m�����"�^L�酄�.t�D_8;�J�A3���B��P(�`����v��ˢA�m9���0�~�!����k׮͛6mڔݻw�O�R~����벻v��!��G�ꩧ~�l�X���.������ӧ�������ϊ˪G���D9�tӴ.�s�hoC���u�PXds�%n���*�@L�N����_8j��Osy�����.�|���SN$� 8��:�U&t%ԩS��������铓� H��}��U��4��tu�ϸ[@<�ςɔ@�&�5����!~�# ���ԶT�U5�:1�� -��a\�8�r�C����q�G���cRB�b:�΄���`�����者��^�7 ���y��alO�6�ұ6�6V|�x � ��	��p��g�EeE������׿*"��	�N�	eHS�t�X!#��H�A�-xX�TL��Kz��%=zv���J��p"�X�̀�ѡ��[�g� nD�âp�K3 �I����\�U���[��t�� �����k6��Eoɦ͵���M���x�
%J���D�lݩC�RP�'T!�Ν;�����#+��\;�cL�#������c�Np��8wd���C�5��)`)�c���� �G�M0�[Ʈ�y�|0>�Đ!�Ǌ{jm2�X͎y0O����FW�Q{�JZkF�SV�SZ�L�c��Z���bi�D";c������7���l����xx�c������q�Ԧ�ƋQ��:�?8���$�?~�e߷�5bY[[[�]w�~���9}�ر���XU^y���|-WE}r踡��m�}W�c���-m������tH�b��֐����;W�t�9��<��%K*���;ӦyJ(����k��*/Z���JE����r�7^1p�����������nO�-�C-���Z���P�:D�9 a �K�R�����xD��b����`(2ð�R�B��U��n�/�H�A���D���4�s`��&�3��1
�X��"��[o��2x�p���ٱ�t��ݱ��8G�  ���T�S�A�g$�;~'��v��t�S�dG�Ƃ�F�8��ATU"�����^�]�!n%�e:#Z:�J���oS�����uIiI�D!q;�R��0
%�h���|Q����G��}�H�.����L�l�:v��Y)̕3`�F���&��k� �~ю�������|�� t�p|��<�ثT�Z+��D8)-�D���r��������D�"%eU�i�v���z\9�!z k�����vd�4Xi?�#�߀��?��rv�#}8��k� ���և�+��6�/0v�p�������b� j�P�D��NV�U��)�����G@�3E;�ҢY�������t0Id̬Vk�b�4�in�;=k��|o����C�wo�6hP�}zr-T�5�_{����H�L,0����y�6���C;��+��~�}��q��Z}�G١S�N����{

�����(���=�bݱ���FS�$P��a���!���[C�:�9{���n}%ׇiŊwK���9i3}z"�p��p"�5�H��d2���^�:u�#F���j�,���3\N�OS)�@י�t�;8U��U1��ˣ�������`pe*�z7�����gWQQ�Xw���D"[�n����٫W�a-͍��$G�(�� JL&BbBBE�D��a�ᄤ� ��R	H�.��ܨNaE{:K)U<�$f<���:�����J30T��:P�J+����E"��1�/�w��9ڝ� &�'��ƞ`~��#A�СC�3 ����5՝���E\��!��.�n��W�#����<@�!��|�H�_7 -��
YZu�,�k�;�\K��蔷3�JlW�sYJ�����
�Q"U]��h�"����&y���使.��j�%i:��T�t��[v��6 P	1�I� =�:�"�-�烎� 2���;��d�t�>���`�x�rh�=� ��^� �q^1.5/t��y@;�I呟���%t\�=�9�9�yD{]�U��3��;M[�������E��]p/���5ý�B�@$i���+))^ZVV��k׮_u�ڵ�G���
o(�r�7N�߽�\����}�Y�Cb�r ��T�aÆ���_�v}�zu�ǟ��p�~�#�aaa��%���Ó�1g�����ؼ屢@h���,�pHl6������-�m��ٿ�<�!�on�Fk׮-�=���T��4�Lh	8�T*e�����N�z��Q��j�`�q��9�[o��l�S)$��!3�-��f\��G��r���644,u:�K*++߆)`���m��.���y���X��Y�|y�/���5���{4�0�=ʕ�������sNi
�VTS�Ǖ��pA휝^�!@$L�p!$��50gK�)bqf�H2a�-:��f�\���L�,�/~�s!	90'dE�DG��d���a�6��<����yO�;��Tרb��D�H"�:�����O�����>lZL�(8�y�cSW� �[��� Z���(�(6�.� �_�zF��VK鰭cL� !X�|����]�d��KZ%�tH��ݤ�I'j�Ie�:�����O�?�=���jf�rǞQ�s�<3�ߙo��z�9�9���wd@	��W��,Qݯ�.�I��D_8K�g��y��
���p��x�w���&1dC�?�|�3���=D.�j���U2�L2n�h    IDAT:ޑ�ĘgX3�N7�ҩ�b��ӹ�����C=tˑGY�}�{��wKo�u댺�]��Z����gCR�y*(��D���y����8˿s�o�Gz�Vo�g܈#���e�

��ry�2P�d/�r�+,����g��Z�[$
�=�PDz���������X��� ��:sj"�%�P�Y��D���/�䒟�q�[��Z?��s��{�a�O�����I4�xok�5xf#4
zccc4��ihn�SUU�~���)�O�^�r��?����I�RA�����W�|�D^�$`P�"[U� ��?�|{|0=ó3�Q����w�"�l^� �	D�R7�l��/i��J W���CcL��i�d|���Ϩ�)QRB���H �^�N���kCwTÚ4�n��*�U�u/�ݻ7�˕�#��>}{JEe��G��G�ax�g$t�T�gy��u_?��o3�LG�;%p�	d$r�nϼ���8�/	egGJkCH^]����қMX$�*@�b
��8(�r�T6p�	/[�Ljj:��(��ƺtq��NZ�s'd�F��� #�}�M���S�ȩѡ��@�~Yp�ca��^�̆�k�����3�Lan�Q��A�Pm��R�48�f, q���}`0':�R+�gf��4I`*����d2�lmll�)��������AMM�������.�7� ���s���3����~Ӊ��q_�B=�!C�<b��[m�߭�i�����?�u��4t�К�=��y޼ǋK+.7c�kZr��^z���e�)�O�6�X�A��%�pD-!i5��F��ٱ�?��_Wy�w��~_�~���fM��b׈HT�x���6��if�������]r�%��0��ɔ)Wݶe���p�����6� �p��ǫP�P(l��r��^�mBZ&L��y��M�TUT��������xW��б�w!T�t*��mJ��"*��jo��>�"�$����%rd�,A!G �T��NOo}Fj\C�#�C_�;�,�2t�C;���U���@8�ʇ�7�(}M�{��*/���Գ�Q�Oz�5(I�ňK�>��q�t��˰a�����W�|�te܆]Ǘ��z�i�3�������jo͠�=1��$���A5�T�II�BJ�n�z彥�c�>-�ER	�t��]�aY�|��7Wz*�� �@z��v�Cǎ��>�7f����b�G�(�=������l�ó��ɨ1Z��1p.(A����ׁq�*ǵ���Y��&0{�_Ŝ57+����u񢌴�����Ί2C�f{a�Q�NB;LB�ΤO���/�C�l������|9���s����n����jCQA��Ҋҷzuﺪ{�~�Y��ޠ���m�m�����e��T��i�=�h,���QG_w��G�D=�7��?��>�����ݧ��#�8\vǦ�����v�'�L�����]�3@߰tqٖ7>��$9�hlr�ZZ����P�ڤ5)����G���	}������������f�a�B*����*5 z&��ѣG�����?���]�����>{��NOL%�|M�
ȵ��M��<�㐍-�����}3��x�7�^3��u�Y?!�13�N���	9 ���k@��AB5j�*!��2��Q�L�L�9��ę^� ���
������{,�õ$� ��#�x /^ rh�92���Q������ A�1;�V�ŸT��om�w��J�̓O[*���'��@�1qH�Q�ұD������I�_�����}�)bU�2^�X+D!��%��1��A�pV��;��ȵ��ȵǻ��~�K(P��Y|�~�F���?��]͒N٥C5$���\�R��)�p<� �0��'";m���f�
���?�ol��D���p�ْN��[�Z�)���3�=�4���V�Ҿa�F|�9�٢s(�s�9�s��!
}1����6x)�v���g�3B�{&�@�ߘC�f)摀�!�=C(q��HP͓��X��d?������h}(Z��y�VUU->���u�;wF��.98���{B���0l�� }A�"���ng����ѓO�������oAR���;��~z�,�����;��������U��8�0�{U���#[��E�]Y��Ԭ�/L����&N�[�Ѹ�6�1�H��ܯt��_���w`VUW�߷O�C� ���b��&j�����KP��Q�(vE�j�$��4
��QA�N�;�����}�Ío�2���rxxf��sv?���Z�:�g��V��O�;�ޙ�f�Hra1���� �
�V�;�ԙ3g>�Y&��s��}��?ޔJ'$�ӆ�ʝ4_SSmN9���<ϫ�e�C��:�e�5kV�7�x�,��w���)�@@�i��Ջ�o��eͳDS�G��0�mc�sakA^J�̬NPq�Z`����;3�c�r����w���'0f19�g|����#��>����(�KQ
�/���H��XAY�����a
��=���lqI�%�h�A�d��}13���k���C6��X�h�ޠ��(1Cw�v�	.��G=����u>C��;ω�:�|�9�|������,h�xBf͚&s�-���>��2�ڞu&M�w�y�&`��ј��Xߺ�-Β,50"�-?�A I���r��d���š�-��r.H���]!eb��v����"m(�Q�qV��Lߜ@��!�0v·�N�¹���1�Х��w� `׊��޳�o�	��i���\�����c]-Y'�𻀉mmm�T:ݘ�dV������_�zۭ���#6�3��ͻ_����=���O���|>�p/6�� `�LWUUD3����׌a�Gw���M���<������>��ˮ�׸�~����n�~߱~�ӝ�K�2��z��E��������Jڣ=�7P���Ǚ5���)�6M���}Ǝ�4n��]^����-������-a^0P��0xM ��l�ͮ��kn�ѣG���.��ۿ��{w���a���EǇ����w�}��z}}��EEŗ4`^g�_�`��׿���Ғ��t�6g�s���bfD���A ������#�<��bN���X;�DL!lB����`i�vX{�!�W���c�w�F�1W��0�K����ς���
`�p%�����=̯앟���*/.΅a�>�������|�!���xak�dҭf�]�1�m���|H_SP2� �������Oe��H6��7�7����$�=�qX���iqik�w�l�ѻT�1�k7Tek��kg�f�X���cY*,3�X�ZcA�qH%Җ�����6�rnm`B�$d� (a�sC�>)���������qI���^)-��w�AY�`�rpv$�)�?�\\~�DA�Kh$ &B��<#K ��H���9Xs��h��X2f���.�~ �J��M����e���ю�u'�	���0O�R��d������7��v\��{|��n����x���pxg�
��L�С1���m�t��<~֠A#�,�ڿÐ;��j�_^���C��f��v4�P�t��y6(>�33�uCg�����֬���=:(�n�1Q������bZ�iS��_�����u��X��Ɯ9�z饅��e��.9��
��z�������1c�e[n��&��f��s�:��+W\����S��CǗ���ӟ�"����-�,�����;=sތ_�r��k�̉D#[�y� Ƙ�!
Fe����q��Y��Xa��<�];�$��Br�1Z�7�D�*��f��--���n��{"A��p��='�u���U�q��X�R"μ!xr7�d�^9T��ؤC�SeAa��q�/�%W�5��Y=�h6�E���#̨QC̀�=M�j�E6}k6��8�q�^���6�|��o7j�Ҿ�z�y�z˅���]��C�1����S�x�+!��Q��ˮ�=�	����~C�e^�x��܌ǆT��Y7�D�-�X�xŤ�9�e$�n��3��h�}|�%W�4o�^HtƢ�RW2�S��۔�@ I΂�~*[}���:�.,�(�gW�&iʌ[�k>��<.CZ?�ؼ
~����r#�s7�s!s����%hӞ\\�ao�$8���*���3MMM�%��K����Ço;w�ԝVx<������z�UWz�'�'�)����XU]av�i'@����WrȾ���}�sޯ]�y��n���C��{���[��ٳW��x&�|!����x�R���;w�,������=��U����ʹ�S�1�]�����=�>��]�x��}�=��}�`p�����U��f������Ϙ1�Q�Fm����>���K/iin=���Q3���T�L�L����v?kȐ!�wE(��w߾Ţ�����v��hTW�XbQ�H�G,�Nqi�-��駟����7�x���������<J&���L��'aG�f�S@(��uB�R��c�"��- �|��1*�Z��+��w����!+��+?��|`�0���F[�M�]��Q}�3���R�6��ʠ���f��[���+lzP���Rs���H[`z.��RW�Z&�;��\�@pb0�mk��Zϥ1���+֙K��0�MSQ^k��ܼ��+�=�hz�Az]���>�¾˕���u��s9��N&d>g���8!�9J�ʞ(�IL���dU�a8�+���X_1t	��oϘ#�q��=U���X88�#�Y}3c�<��k�VL���e��O��w��.�4������ i�Ri��Z�v.r�/S=�W\� y���������d��Ҳ�;��#^�a�6Ya�&L}���C�}�yƘaz�'+`l����PC<�∣~tWU���}R����Ew<��1_�^q�СC�f�u�I�t��������B=]�������ly��KÑq�Ƅ#�6��#�9�0�)_}���{�|��u���)��G�lѢE�gϾ��` 0����R����\,�Sg�u�	t�&��?��ÞW���u�d��t:��g�EAb6>ycL[��ź�6�ZWW��7yI��3s����k�ܝH$v��	�ۣ��� �ʐ&�D�D(+!�?1�=��s6����|�z9�Й'�E	D\�U�T��� ڴ�%��{� �G���Kq��32�ӷ T�/��Y�2a�
��9� ���̺�r �dh�k֬���47��2�U��e}��$d�&*Ș��8���(SZB�:)^a���nS��R��CS��,o_WC���1�cp��cr?S�w�]��q�Z���|�i[C����_^x�\�m&7������l�Y���vϢq�ϼ0T`ӪU��0J��4k㓹;ߏ,��4y�{��%�������+��2�����9+������a-�\�юD40M�g��_m�<�?U�C�$䎶8��%��W%�!Y��rY����ɹPM�Q�f�U���*�%_�����u�q�^���&���E�p�'�wqqa<�N/�d�������s�!ߺ9��3����Ez}�z�X[��,���2����1�N�{�?z��w��������|��'�����g���8g~�����ǅ]m�ե}�3��Z���_V�ۏ��7xZ�;̣�涨iO��A��O8���G�eQX�O?}���W_��x� U*<T�r��7L�����?fҤI�7q}�K�>���sf߆a_��/gN#�u�&�8���[��������G�.y��oΠ�^��h$�D`�F�y��x��p�������Xl�
���a���Τ�P�|�.�
რCp���\=����2�'h��ړ�(A�̏
wc<{^�0�3N�2�ў�鞰34瀱!h(�J��_�� ��3�i;&�Mfm��l2j��כI5���������>�6n��e�Y����ژō��9 ��aM��?n�v�����3.�
��7-�"��&�H����y����G�5�L����(�n��#NRT�4&L�0,΋��r��(P{���D?����la��B���J��Eg�1ʬݧ|7�r!�<gA�)mX�bNg�|&s/�����a�|���^p?�5���PȄ�˴�V8��U�E�����3��\���WR�@�5�I�%Y�=��"-���ʊ�w����764�{�!�޶���k�3������{7����1~�`���������7��r�qS^�T���<ec�ϛ���kW�3j������z��������3�٥���^�\��秖�E�66W��,��@�D�4��ļ�B����i�~����d._] ���_�%���I�@ d��\a��Xtc�;p�1^��Ec���?��_�i�ቬ}1��L �{�Ǌ��KG�0����%��C=4�?=~W*�r~<@b|ʀ���q��ɝ%*�Z^x��oC�-�H-��%w�w��B�0�s��`+��1�����	Ҧ�ˏOg.��$�@�����B�s����,Y�+^C�� W�����O?]n��ՙh�dnueҡ����ihZe~���f�q������p{-fn3ʘlGA����}������EZ26#(j'��;-=m��������5ff\}��p�r�).Ҟ4i���_�VI� �@��`�'V&��B�B�����7�A�!X���,cb��py���k���'2Ë�ڔ��}��-+�Ί e:�I��/μ@eN�SZ>���<`��}���j|߁#�1t���(�R�:�@����>z�笟�%K�A�������� r%&� 놕�������/B�»8�����O�(_��0���9��?��t:]�X��޵�ö0�첋Y�v��e��z葋;�������[o�,^���u��4r�m�C�n}_mm�G�Qե=�曁�}�����k��&����hGMk{ʴ��l5�#f�jQW.�g�}V0g��W|��šP��?Ow�}�r���3�뮻�M���>��瞺+���J[0t.:�f��>��2hд!C�>��������m�~�ٻ|>߶b�̕�U�����<o��d�Д�oQm�R����ef�Y8:B��hm
mY�l}@"[�i_Ҷ��D�G��@P����Ah!��	��V�sI��9�(~;V~��J�ÏN��.�-c ��:?��8�ma�c�V3h@ws���LYY���̓�=�4P�XF9��v��]�RC��s �.��#��c�0zy1t��� ���1�P�y�����ko6�MQ��74Y��
�d��d��0�LƮ=�W�&m�`�0��T�'�Y�%K���e}�~�9����%�%%`:		��m	��-�=L��3�$߸�9}ӯ ��=��m�8T=�!���r#��%����WW�����5O\FUB�;���`�{v<.�����Ug�p�L}Æ��
�8��5/���W��2 \�,h̋�����ē�v���W'�x�o�n&�oB�(��1�����x<^&���	cw�ѐ�|駟,�߳n���ץJ�7�æ>C���\
��َ�b��x�2t���׎)n
��k�\���qSRXd2^�e�--Q.}��v��9�����~�h]����>x��{


�Hijn�4/��G�����9s��[���\��ox͝;��3O?qGKK�0�Y�X�c�|�gii�9��n��������o�Ϳ|좋.:h���7f3�:BCHh�K$Թ��7j�4A%l�!�!գe-^�ؚ\囆@���d�A�BxQ�6ڃ1�Q�yғ�Z��m�q��l�&���g��P¨<�0t���F�E���0Nϒ�� � 0@0� `�̹{�ٺ@$'R��W����>L�Jo3W\u��߿w���8͙ح�lG�����1t;qWE�2/�gwھ��ؽ�62����!�Y�̯!s��ߙ����),�2�Ma�5!�f�5�;�W<�kKn���Ֆ����3�T���`T郉qv��X[�|�sx�\�6ڀ��"����c�dRȜ֎�J�c���&��#A@~ga>�W}	(G{��`�ֺ��1/�@.ɋS��<��U    IDAT,1��eHt��{�U��W���Γ�6�H�I����@9`<���X�������?d�`=�{�RX��ј͵{��@a��p۫�G��z�i���ٙ˾z��P�?��+c��Q�h��q�2� ���16,rɒ���v��]Q$�_���]��ߞ;w��wޞ�#��3���d�m�����
Ms��Dڢ�!�ٰ�4t��w����4h����ܲ�����כ�	&\�-�}�_���|���/�p�ȑ�V ��ν����ǅ��^�CE~�<4jԨ�����aW����{�r��;.�x�'�Ñ���F�y���Ң*LF��$&ĈD"h(�$?<ē���A�sh~g�~^X�}�|�����B��Ч4m���	A��G�K���81��N.i�%��#r?�Aܸ�W�{���\aQh��R�s2�2������x��3a�����дG�-xL�n�''�Q���D�՝Wh�K�����󋭸j��yNkg=~��8$�&�M>��,�������\����?6�L�4��M*㳡j�H̺t��\��nU5v�ڣa���	P��s֘�?~�y��7���ϫ<�1�Xq�G�U&A�&���Z��N����Źa�Ĥ������"!���_.�"3Ĵ�#Yy�Qh�@�E���3�$���w=��G�SEk��XCEY�����w����fpr��UD��Eii�{���d�k��c�Ʀ�n�l�&�J�Eb���d�d2Y���Zd��)����7��k[{�il�q�=�L>z�1G�|��^�4Hm>��#�n������A�L����G�w
S�o_|��;�qɰa��2]����.g��<6��ʗ^��W��Ի�� ��f�CA�Le�ݴ��5��E��v��!�F{l��r}�����Ǉ�(*,܇����l_����X,��9��S�v�a��G���>�����~��&{���G�)�T�\�/~������ݮ8 ��?o��//����h\�f���o������̎�#C[�u�]-A�t*`��|�<���� !��'�=�Bpif�@�o:�si�`���e��9��|�Ҕ�
��%B��}B@��C "i���
kb�b�h�n�xy4n�l3):+, ;^��E��С̩S'����M23�`�d,0+e
Bŉ[Өc֮Z���w���}��Y�l�9�s>y�a�i^����>�,h��J�-4�y�̾�N���n2ig9oc�3�*"-6��fD��=�F�`��r��4����������7�鰄(�\�q	f�+S ��ș�/�:��~�\�L��a�����
3�+Jr�}�_�8�2�s?{���;K?���Fp�X�5��5�����.32���l���3M�M�]bs�WUu���tu"�D���ݬ߀����;ߤ��2��R_4������֭���7o�PK����Q����֬)�]ĺ����י���d������=jk.?��S��իW���f]�̙�����3'�L��؇�+��^`�@��ݫWf����l�Î�<x�������mv9C_�hQ��O<rz��95��\�hh2!L��.l[s�iNg��`���cv8y��i��,�g������|�Wc��Ǔ��k��A	]�j�
���z��~�Yg}�)�������U0����(����不�z��l�ͳ�g�s�珗�4�gϞ�z��K��l�����l^��WX��-b������c6|���A�*�a�YOb��9B�7Z�����e"G�s�_�����
sb�BC�eZT?�O����f%��)$f�8埔��M?Jj�a�G�8_�ʤM2�4o��9G����2~_�Dc�f���́?��Dc��}���Kx\�))����2�\����r�K �az�����`I� �~�1�Dʄ[�f��כ�� _{�ik��p�5������qg��Y�îE,�P�|�.'�,f���{�m�6��w_ff#����8��?!T��]�t��ٍ=�}�O��|��K �~�W?}+�� n
M�oL�[m��.8�|C�*��ёX�@p�	cD��ʞsW*2��s���M��"�lv٠�C�����6��aÆ9��?��	��i��h�G[�����J���-[��_���+?���A�A*��|�lsK�s�&O<y�}�I4���/���'�t_6���
�y:�x�A��������;�����1��?��]�г��Z���"��[�}�k7O2i
�
M<�6�H�4$����/4��?�uV�f�[�zu�UW]>��=|~qQi��`.�"�f͗�E�d2��3f���_���.�W�衇��;�������/^~��l*�o7nܜI�&]]RRҩ�{��z��,��?Uwkoo��n�XJ뢞�Bv����a�w�ٓ��he���ߡ��)�4̓�B�a����&�cf�_�o�3� K�PXڸ�b�ṶB`��(\f�יּ�XM3�W\1δ!_$���>�:����hĠc*MfҦ0�B���*+JLmM�ii�7��u7��~���3YWJ�{6��ׁ��A~��X�y.�+߯������$��k��i�����������M$�b�J*�C�=d|`�I�0��ͺ�M&�ʚ`�ȤA��ʑ�Į}"i����
����YSΉ��(��\&��z���P�����]���
Ӕy[a�x�MdD2��;L��E���~�7�����pf���O�s�W)/���s���9e,�$(�'ᛘ��z뭎,v�zF�u�����;�]�90
�'�1�E.�rР~v,�����D��ƌy����ª��=���kG����;�_y�1����/W�|�g�҆�#�XAޕ7n����z���M�4���4��?��'�x����}�^c���d�������x,qΘ�vz�����M�!���]��ȋ�ݸ���9������&kc�!j�ēYS�1a�oU���q'�}G�=����N��7���w�l�ʻ{����O,!.+s�-m�2%��۷���կ��T`܂��1��Ym�g2/D�؆fy�	�����'���{���������͝��--͇WIÕ���.fW�8��l��L���nV+�dQ���*���0Ee��e� �g��A��pҧ���jf�����!���l�Ҷ6+lж�����=��� ���0�&�s�4'�� .��OB���	��?��ck������3�t��A�Ǔ��e�IS׻�	ѸZ�v�����?�dR��� �`���5��"w������k��ߦ���=���� ��q�x��C�'�ͱ�j{����ۯ�in����5&,2�ᨭN�ZQa�I�3&��Z���d������̽^�cq��N~g�X���O?�<��{!���	"�q�V"�v�,�ݓ]��О�ɹQb�9���
ٍ&� �R�gd�W�&�_8�g\�'�hF�����[-�6���C��"�u��\x ��,�N�3���.-*�~X�P�Zֽ����O�zۗ8���M��/~��G[�44���4qٲe5:�����0�K�x8UZR:��'�����l������7�̜1�U_��U6���Y�����#F|����+���Ip���$�)k������ߛ?w���޻�&�=0�v����=��L"eL}K�iO{Zc%e����/|�a]�7����.Z��}uu}G�Z�ږrU�$4v6�m+**�{��W_���8W>��s�������C�>��K��L&#���{�
�L�f�m69�!�{��Y[[ۤD"QG8�\�(d��IQfwVZi;!�\h��.?�B��b��3W��}@L��UZ6�B�X��`z�g�s��]�W}�E	�!���0f�̝U%%�Q��/t3{��`he��@Km��s�ޣ�
��T�dS�@�g}֍QVZhj��L �����gv�c�m�cAL�J�v0�f����i�.�iǕQw��e�������[M��ܤ�1�#�κz3c�L����d�k��c��5j���LgM �p��w�@�^�-�L�j����%cQ����
�--f�ȑv�^y啎�}����=��u�yT�8�`Bk{���X8]���L���9i��#�]L���.��(�+�z>�S�Z��QӀ����#�
P�p�JU[�o��9�̃�+�,�Z��\Ŧ��쥞�zM/.�zc�w�d#����zjл���_~��hcL����BR�z�@��Z+�;Gyı��P�g�$d�.8�����L&Se��%�a}Ǝk����>�VSy��{��%���DF�Yc�V��瞫���O_���?.��� ��j���T����֨i'ӑ`𹚱#O�c��.��p ��ν�ʊ����e���X"��x<OM�2�I�6���i�����775�X�>3`%$xu8n<x��{�׬��nyMM��~�)�<;`��G'�X��l6;@L��9������N�y��5��0ċ��lC�$���Bؤ��\l�/����b`�BCd��@0Y]�*��cA���gX;�:m��O@$��#�W1ڃ�K�ȼ
�f�h
S1�)�-�Deu��޽�J���
����L:n��KLUe�������'��ۍ4�t��D3�����1�U�s�g�����,�<�٬�A.�����|�Ҥ
mj�D4nM� ׯ��*��R��k����h�Ɍ͜�He��ﳡ��DIK��䥦[~c�ǔY%���<s���B0b��_΂2�_�oΐ�Gu�s�)7�ΰ4\�� ��s�'_Eu�̭�?�@�s�l������=̃�Wn�#�s0c�݄��{e����Z\��
i\B�+/<�ཊ��l�S���_�������c.?��N/�4w���/.X03���
�V�P�%�
���5��4f��S�8w����%��v��s��^y�WŢ��f��""-r���Ͼ��kC�����=bĈ�:���Z�Vzë�����~���ȳ�����lL��H�i�L�)���������:���L?�n���^���T2S ���:Z&��5o��>�O����dO>9����̻$�Olii��;!n�X�2A�Rz,k...~}РA��߿�;555M�t:YTT�...N�B�L0L�p--Me�ي�������/�\_��/y��'�"�]��lOe��0��(�j�9��V#˅�I���̺ "��D@Y�xf�BD�s�n!�\hs�\��0�blg��e�^;�W�1�R�3'eSH�J��C��D.5�1��w�������h�hfX�� P��޷o�	@��z�����p[�	<�W�����5��$h�>�p���cL6�>ug^�i�b�0rk3'�[Τ���7�O��:�F�MC��@Ҡ�Hk��w���6|���{����W_7ᶨIe��=7�p�#��	��mHc��CT��[���$�]*I�q��ʎ:�6�:��\fx@m��Ť�i�'{�z+1�	O�����w��{!�l��MMV�S8%�s�/�O�������\F��*�
��{�BU�����sR��#��!f0t��A���?�{�uɋd�W��S�8���Ь^�ʂ��ᦰ��m����f����ܶdɒ�Gy����l:3�
*����Y�d*�Е*))��y����^�z�w&+|���n�����~���n�Wَw�����L&�ط߀S��b�����^�o��3��g\�_�����xl@fC��D"&�Y��qo���dfu[���=�g�v�c�����g�wnįtל9��\���Ҋn0t��җ
A��'>��VS����7�?={���]�ní�֭�"1�������?5�N�7x��������I	����~�?��f>�'
��` ��$�H�$i�M%S�@O�7`��E�`��6���`�'�HK�$�w1��P�%>|���������qˏ�'������KK?�;�*F�5Q\�����k��`.00ƨԙ��,�kʘ3�p����L�<K��I����n��abG `��ý4�?_f5��*�lV1��e*����6������T�7mB>S򛣏>����&o�a�T��U�ܾ���I��
������	9���S��EٌK�����h{�W��+�4w�u�y��7lvkn�S��� t�����kom#ď���Ja�w$�ٳ��YU�o�ٛ5��F���x�n��{�0B�V�!
��Q�??i�3�x�K�H��v�m�_��G� �q��^���\�,��<��ιAh`���0�9��3�4s�ε�s�p0?%�a<�m�X������1W9mqn9w�@��=�f��߿������6��5�o�}�}��s׮]7)VUu�g�uC�iq��ǧ�~�#G���3�ڸꪫ=���$��텛!�!k�~��+*���_�5�����Nw�\�S����Kw�Ѿ��۫����M���%a�h���Mc4��RU�Į;��a�ui��k��v�W_]xo]�[��C`(�l0�h,�ԻO�;/���+��z�M�p H�r�g�ѣ���U�V�@``�����Bܙ�C�>���D:�Ng|~O&�N{�'���b��"i��>��D4?�=p�������y���H��E;E;�1���L�2�)�WhZ��0&�`=��&�P"�S*X���%�P{�8f%b�D����g͜�X���>Yw�_ *��t48́��{�ˢ��	S^Ui�ʝ)�;a��755���f��������I��n�f�]w1?9�`��$L��e��)���9�ݢ��ĕ�m�U�����d�#լe$�"�ɐS i���BC�^�ļ���f���5K?���|!�L�L{4iZ��&��������g��'H��EE�w����}++���b.1]Ʀlh0k��~�� ��w�� ��rYS.�'���9�{�w�~�����L�B���O?m��1+ԑ�s?�
�~�A�6�+gM`� �m�t�M�Y����/wX��N(�d��yK��;�f~
�{�����鱲g��Sv�)�P�[pD'q�l6��͜��䓏n��[�P��e����1�&7aҞ{��q'uk�9���F���ߦR�j7T��
�ĉ�g�]�����X^^ץ�7;sn�)m}k�ӧ�X���o��d,hi�e���������I5�LC$j
/��c�Sv���M6s��E�?~�{�{������~]}G�F�T>���I����q�'�0aNA}Ιss�{�y�Қ��� ��hf%��v[bՕZ�������,����㖹O���E`�&/1��h���C�o��aԘ2�I��B@�C��G�v��	�$m�ghGfM�ЕVk�y�0k�V�U1d��mn�\A��e>|&�jq��a ܯ�t7�I!�<�Կ��Z"E���0�t�'v�H	���;�I$l�o46A?��E�g�n&��b���;lg���������l:i�I���qXQ\�����Xk<�U"1��E&kO�P!)D&����3�X�<���ǟ6k�4����ٰ���dO%�.�\��2���b�Ѱ��Օ��;-��g�8��r$ ���,q��!g	7��b���$P"�͜9��q����G��g$|�j��bl�w�y����:׌MEY�:��|I��,H�=�i���K��|��f�w��q��`�쿘v�<�9���U{�z�
y�o?z�)�&M�sW2��_|������|媕�!�B ���.//{ﰟ�t�{�������u��?[vE:����_X� �(	?��O��\��C���p%��{��+�1��ŋ�����5�䔢�HY���d�1�Y Q�=a��f��,��}�a���g��Ne��k��V=k��WV�W�D�!p�l��x�"����{�#�_9��{U�ō�wƖ����˺u�����K`
y�Q���x��|��j}�9��K�r��bL-b��k�8�{!rҶE�e�'}*ޖ��mHV��@��
pG�B���2W��|�M4`��o�\��3�ỔT`$�~��yU�� d�w�q22}��dX{���{%�a�     IDAT�Ҷ�1"0o��s��_�n�P�`�\�oΗ
���%1[Ǡ[u�A��J�M���f�]Ƙ=������i2I�ZGr�_� 	��.��lh;@�:�t�X�/4�@�i��7�����f�����2�7��ih��1�z��4a��\~�H�:��x����.uku�ӬA��6Z/�a��[z��ϯt� ]�\$�I����p���}
3c]y��t�<+�����kf̘����q.�\�.�e}��P�	��)p$k���_�=�/8�>�I��9��|j�s$���U'�ɐ�'�>�3ڴ��]w���O<��΢5���k����?���f��G��d��	Wh�����=�w�a��Jg�c��/���_��m��t�u��0r&w�xᩩ��8*�8v�������W�[c蠯�����׭��,����d�6���L*�4����Ϥ�J�����	3{��e�k�2�8c���������hm��eU�8�%�̼_4��Ky�o;3���ɓG�чg�����d*!8��x�U�K��ܤ}Z���u�6�ST:@RB�K�r�5��2�)�bÜe�M�c�Y�F�h�f��Y7�目�ǭx^�T��|���q�@����Ye��F���!�<�ߊ��y��p1xߣ�+,�~v�X$�M2W��.����
_�go���Y�C�5¹�˘�ZLyE��ի�!k21o�t�VmF�nv;�l��`�/�T<j���dL:��YkhF�J�M�����c��ini7o���y���/3�`���R&�Șh"i�Z#Ĥ[kD������9D3��̌�0���2SY���F�̛�a�4��ف�]7�J���B����GֵC;�{�^p��8c_"��������v �i�J!��I!n�-���}�>�'��?�ŝ�PGl<�w�?�09��HC��.l���2�8@Xb�Z��l���s�9�����av���p�˷'���#8��׬�BPEE��-�lq�	�����&Œ���n�=��&k~��a]H���	3ĝֽ{��UU�&n��v]���Y���o���o=�Ј��{GY42������M���C&��GM}*�m
����}�n{�K�rgμb���~yy�p���̅�p�s�[�����_8�����τ	�}��g?�d�?������Ge!82��S�C�QB����:��G�v��ᱵ�s�]�ǎF�|x|�s��1$>�r�;q���
$��!s)S�H��^D���|��I
A� ���=z��.bO�]���8� �@h�c�{_/�D�&�N�z��0��:��9ry�?J�J���f	zJ̦Ѭ��`	�e�%����#v����f�N�PaQ��ӣ�d�K��1�ӳg�<�����m`���$� L���|��hR��J�����5�&c ��L��3�τ�"��d>���*h�
�I?�gn���E��=H��\B��^\\n� Eť��`y��Zqv9��2��}a�re9E��3#�p.��x��'-�w�)Ab",9샢!�G�'�`��ɖ�"8�Lܼ�|�q��+w���M��5�B#?�����ӭ �����[;��*�\鬰�r.p!��8�5u�3�ø�/��TVU]s�)����|��<p���>7� T���������m����{��;���O�r�WN�r��zl��m��`
�B�]5j��z���������w)��3��R[�*C_��K����W��c��#�����MQ�!�[�qS��&�����C/���w��?��{��|�D"�h�C.��P�r�1o��N<����O�4�ג%�/--ټ�����i`he.��Lv1[�3�W�Xm��v(�|�� F���8mA<�y8����OcB�P�;���}h_�1
�+ӻ4�c�)�I[����9��>er׳�H�D0
���8ũ#���)K����F�6�gy���92n��Ȉ�k>��~��w-C�EeZ¹җ�����n�]��1��d�
6K^�IƩʛ1�lڔ�����2�t&�|��[�x�w֊>e��X��z[�-� � .�1�X�d3>���p4f9��V8�8���)k���������u$������tj:��������	\I��ab����Cҫ*<R�\� �=�i[V)��X#b����?���@���+��,#�ߚ�ss�҂p��@X�e�]f]#$+���oא�΂��G��+֜�q&�W&}8�ejc��ɬ~rؑ?1bD���Z:��ه���k7��U�׻�����j�a�**�~|��79�ݤc'�t�'7�R�:��,�%�k�p�-���;v���}31�[e��,)]��}'���/*�F��k�M0�1%�b�7:������i�h���7����KKƍ����7̚5�����d2Y��FO�$�f�"�Ȧ&]��V�/�sל�:;��v�7�=��c�[�~TRVv`A(ԫ���L&=�I9B�|�b�wQ&5
�U	m�#�Zs�#�t�yCh� P
5�Y��YV�B�X�$����1)Q�L���=���yM�� �b�9[�si���6Ee,f�.����hp�/�'�A>���;��iK��@H���[��ȗ�+K��N�>�ӫ�
~�!!�_�Ye�Xe�v�����\]�� ����ծ�M*�L����6��,���1P�s�;����,B!g�a{�6]+Zv{$aⱄ�Ήx �ݏW[@F89�i�{�{��e�Ν�&i8��������1L|��'i��, �0F�Qg)���#M��+B�������-��^�?���S�v�>��Y�`�<��)̎ߕH&߿����q�O��1ϙ���{��&��b*�"ӿ��%�p ��Fa�r�>�+N�=���x~�NcN7n|������1��W�\qF4-`<u��w������4��g�wA�0��K��M=e괶p�I�d�\�_	�Z����+�<�v�e���A����5W�[e��[g��|����CLc��7����uMK�I��=7|��:⌓;5t"}�T�<�5�4_��0���t���L&������_|Θ1c�L�8�S�_y�Q�d�,-)�3���7YS��z2��񀡄
�,�@�0!"�0TWw �`
h�`��[���^�H 8����I_�I&rL�<�D��4<�kL<��0� >RLl���K;a�Q^x��IZ?&f h<�P#��P!�2���������0咗9�v�'ሱ(���C{��G|��b���
���B���NCsV�D���A�Kx#�[�@r������2#Z�=�h�t�jI�}M��Vh#;�9ׅ,P�q�a��Yǰ}���1(^�v��L����0g���R�>Yx��FY�xF@N�g��,I.��Eu��i_�:ڭp"ӦM3�_�߄���5��^}�<n�!��ƬgS�	��e����1�G}ܺ6� `n����Yk�:I8���8��p�\`��]���1�@���w�>{�q�޽{���x��w��殻nI��ai�'f��?~_p
�٫��ɓ;��>5����ϼ���1�R� k���F�j �xȐ-&o����"H|M^���o���������pv?Oho_S�	oh4�L�a�J%L�5b���&,��z�V��q�Ov%@�n��k��.+/��<?.���>��ɓ'5aO�z�M�V��ۯ�_߰{QI�djcLE0,�!J���� �ZDI~t�L�L�\"�B�˜��CEK�生�+��ye"�B �_8��L�̀�#���2�)��%�MJ�Ct��V|>�y���#��E�ث|�:�B(j1@���? iI�����ӆ�L��%�1Hg�5�?c����������DV	d�!��[�P̗�3�|W�+���<��=�+�;}�s��!�������4����r� g�~�-@�Үa沞�=������{2\ �͞�7�K�qc�=aO����[��0t��yb�!��!�?��U��|~�O͘1c����hq#�q��W۟�߿_+b!`|�)\�Z#�0'�a�8�a����0�D��b�˦L��jgӚl6���[�/Y�dV6k�S.�/� �c��=�Y������i�-wh��o���>����tf�9��ڞ�-ChZRR�ҠA��>|x����y|���z�7�_���{%�'�D�����M��͔WV،Tm��&K�V�m�U��t��N��|ߝ�,�����~�-�(-+;.�͖���y��tF���Gb+w�q���=��G6��ڿ{0n�qz�3�-��ok��$��ꪪ**k�u/�p{���kk��8�=Bd����hG����^��v`%1=�sI+��¼e�f]lR�\B��Cg<֬����&�C�y��D�!�7!��.��`!�0~�%H,� �Xw����oiAGgR�pn�u�{���Lh�[ *�Z@�Cb�ik��g��'�"�(U-})���'�X1o�J�S�2�\� Ɔ��N�8w�պ��{]�Z�3m���΀@f�G�
�h�e]�1;YqH�Y�[9����6�C@O15gaHt���/�M,��H��x�q8��Y��ń�9�\�M�=�Q�	#m)��gi��G$ƱGc��=��c��/Z��f�#y��˿�s�~0�|A�a��C�:����p֟tS*���2k�����lm/������=<3�I��o}�{cc�5}����m�9찣;�8�駟���o�u*����<��zY���2=zt`�-����f��7���$�r߷�����k��Ƿ���Z��X�h�,*8
�x8f��	ӜHe|�'���g?ab�Il�ݧL�th[{��7CÂ�)��e��߶G#555�����9r�~��͛W��_�֯_()���٢`kCCͪu�vٰa�N�x|h<���b�>���Ř��:����� ʁ 	/��{ Z0H��#��Z����Z'1*�?^\5�������z'M�x4:���(&�g!�P�LT&n8�K�C P���0?&T�w�1�m�
��we�+m'c����f�8/$AsC˧��~�ELZnYV�6i ���;��~wj�;m���1b��&-�1H0��@EJXcUC��'�2Slƾ��2��lξ����h$lH��\�%s&�wG� �K�^i_�vYp7��￿y衇����uFeya.j;�}�qn	�����1����MHw�-.��Z'����\����|߽ι�&�Ɨ�E~���jY���~t������w��T2�UKW�������n�cR�d����s��1��n��n�r±���9�SB�/^\rѴi���7\�H&�%�*�FMm7k]4h`}�>}�5j���2�o��׏}'��y�m�굷n����׷�Xs�I{I4��ǴF⦡-j��O�F�t�c��6���t�u�W}��E�����1@����ˎ��n��u��N:���c��=��e�|�IŲe�z}�嗻F"��niiMZA�����*�ĕ���e����Ɉs��&s�R��x�T��0��e
VD�	��*���Ѷ��L	M6�d\�h�B�Ld<#[D[��_ 8�:���:	� �'B���[>v��1�*cC����n�)��R���!ӻ̒rgH �3w��K��o���(A���]�Ai��mAm�<���iG�a��M@{�(��i�Ƞ�|��2d���e���[�Vք5�9�e��������m��U� �?ɣ�����w	\J-�g���f���bs�Q&X'>��@h�ԩf��A6ck��@<:�3Gƍp�h�otֵV:�OY�xl��b�(�sJ���כ	��_;v�+��{ߗ���߼)�o�ҥ}�x�#�.���@ �OggKCUU��-�=�v�{���=o����#��A�L��8x�z��i�0����4v�n/y<'-����+�0t��-|౳KZ�g��ǋR���C/�-���5bZ|��puż�E�]�v�Gjo��7Wy=�Ȣ������jK=�ل+�G���K.�䮮�|��{`޼y���nI}}}��k�n��Դ�����L��e�d2��qsG�/Sq�ҚD��B�H�)���~��!�2���K�|z�߹������y�!��	s�Y�A������k���B%5sR�L�2+�DT�Ի�y�%d4��3��O"���Z�� �/�;s��\��	�J��4HŴ�#��I�� �Q]�\�W `���h����q���v/d�A���[4j�^~�!cWp֍v��{�C�$��=���5�^�JfxYSX/��/�\c�%�G���GD B�y��О��2BB����X\x�Q̞��u�Yg�d<af͚eƏo����v��1-R��Js��53ϯO  ��仩Ii)�J������v#��r�!���j[


eee	�������+|Q6����K�z�ͣ>����}>�-��EQ���+�u}��=q�Q�6��b��O�>��瞻/���Ct�wd�-�X�k߾}�:tД#v�o��M`�	C'SтYW�_�fv�>����k
�~W����D��������=}��'t�O��t��Ьk�9~C��C�P�R@Jô��j/������M�v�n��rֽ�}�駋�x㍊�>z��/V���v�D�[����


�p5@\)	�qD�	��ںB��wWHa;2+�N"��LDZ �K��K�������.A�x�L�_g�����[�G�ƪy�v���ܣy�1BH�s8����ϼU3]u��C�s�� ��Nhfb�UƩR�3�3 �'muD.�		|���k�ż�;S�3�3o�#����HD�uT ��_Z�|�Z3��47�C�K�^��[8
�`Md�VX$m+q���9t�K%���Y���ʚ���׿ڶ�W����E��˒��\��K��5d�m�r�9�c��z�<�����O7�]w]��k�a��%C�B/x�dYQ&:֎9I��t*n�-�dQqqǹb=sc[�H$V�B�u>_����6UWW////�������Ń�`��ȟ�z2^�'��S�tɊի.[��Ɔ�mJJJ����Z�����8n�qS�?��E�I�&u����m�x�da��b`O��9y�_��n1b�K�e���9��Զ���b,�3gІ�?�����!|-1>O��3���C����M��0��h�At�)���uYl���ӷZ�l�l6�/DY�d^,4�\�ϒ)S��l��ɯP��?uc����_��tÆ�V��lȚ5�~��z�imm��f�R�LYaa�_D��\���%������r��5!�"��43�����Oq�s4Z2�?.�ʫB`�1�W)��-M	�1!?8��F_�+f	��y �����U�b���Y���OŹ+E,��T�Z����.��Tu8��Yw֗��-�\Z������G;�� ���DC�4)�*����)O��l����Hۧ}��Gam�p�ښ�f,�����UΓ�#�Q�
�H�Z�֓Pȕ���7�3N|ت��|���3e�S�U1q�a�đ@�Uv8��	'L����.{	]���;B%Y'iմ+J���	i��`\*�K��׹時
_�On���T*����EEE�t:����"�D"��S�l��l��L&��d�!c�������y/�`�@�������h��'�l�c;������_tљ��-����*�s�U�;�o@_p'���8w�v�����zS���1��ŋ���c�%���J��X��x�F|�/dbɔ��V�IE�����#.���6e����'�|�f������<"�A��7�n W@����ꞙ3g^�}�&��̘1�⣏ީY��qX,�)On���>�l��B�C\�:@�!x0�]v��jD�W(N�)/��KMJ��ӏB��Laz1f��B �U�o��!��GF����|�r(�-M��ʜ�j    IDAT�gʳ7�t�хI�>@�'4z����#��^JY
��s)z"'�6�ˊ���[_�K�+3��Ե�����<?Y�J�
#"�����/FĞ�r�����gج��X�|󳘦�#��u��q��H�b��IY����jvr�H�V�9�PT�"<$��!0p�h[>~r�}��V�|����>��c�$����8od��.(��I�P�R�wA��ߞ�x�㾍@GW�HV�R-���:#+������<�V���wD���}��ht�1�}��Qg���n���}��w����N���;� �+Bv�^�$��p��Qv�y�7;������:��ܬY�&?^zs�@h`��դۣ���iMјِ������}w}��矿�_����&R�夓�?���eF0죌d
�œ����(++{��N�t衇.���}��͛7�W___�dɒn�}�ٶ�W��/��7��e2��ED�1*�y�!"0u.i@
���*�#M��` ��o��}�Y��¦؋|�)��L��y��w��a
[.�4�C�y@�����cÌ
������D�+�Qw�eJ츰>о@R|.�Ƙ�6}�U���A>���%������K��m�al�!�Yf�|������U���\V͗�!�([��<WP`�M��{/�I���Esc�bz��?L@m�]B�N�i�{�zh-����uH���s�;�d=�9���3g�Y��[���p��e�:�r�0fa��D�/�wE��=�'7D�[A�	2zg�`�wdy� ��ɊE_�%���p���fk�|�ގ;��d����l����SG����z�ޭe�a��ְ�5fР�O���	�l�M�����i�w��w��?�Ƞ��~fV�¢�5�K4��P:c�%�h��Mc,b��fox��ז���v�u�YÞz��_w��}G=��jA��}�y)
��O2�����f�������Es���+{|��G���ֶ{8�<���|>�@I�r�hI�	XH!W2A��Js��I�yҙ�����$� ��P�>چ�i'�d���'�t2�X>I�F#�  -���Sf\0{ 	�Wa\��7LK����E��ږ��hO1�05��?������#3��8iX!���:�؎�+���Zo�p�v�?�"'����G~X�����4/���B�B�� Yƒ_+�{����6��i C���l�z!`�UH!sf-8?
=e�� о1t���!no�{��}衇Z�˵�^k�h�p֭���wV���p��dR�9��b�K�[H{�dA�i����0.�����q����R<���P�.U�DSs�]/�D��l�͒��M��j��<h�g;���\V.ZYxڌӎX�v����V�$?��=�]�]�+<t��F�s]�>}:%�M���M��)Co|���������E5&�-���dZ�M��b3㙔i�FMC"n"��Ϗ���m{��ot����/���k�(.)9��(^
�)-��/���M?q�W�6r��NM��Us�w۽���˗/_�gٲe�nذa�d2�ekkk��~B�fϞm~��[@�A�%}C�����\x	�Bؤ�1F�:/?�G�s�,�A@iG~�| }cz��+�P	f �0a��iGV�.3�̛�!8�+_��55u����rN�G�Yd�fN�����h��'��?s�kA��U�{1r����:m���{��e�P����62
i��⥅�g�ʀ'f(�?�b}�^��4�|`�L�{���M)si�=d]�d��<pѮ���^���LYS[d�� E�E͟vdn��D�	6��{��ZI F���{ﵧ�C��]΅��V(�B��;r�'gH��N)�&��5�gR��A@��B��0��k�w����������X���l6ijjzk���7�~������v�B��m���z�}�ݳ��Ç`�`̈́�`Ykj9������nw�^{����������}���N:��������:��z����D�o�����kZZ[Mk*e�}�e��^wzڥ7zF��2�������㥟�\QY1@D�]ZVa	��b������ǧ�}����_�����{��/_�ɒ%vI�R[ZZ���Jl.��o��s#߉�K[�YW]��<?��a������C��wW�S;�� f,�;D�{ p0N4w.C&N>Q��}�a
%ӧ�qb<�Q�A�%����E�����
�oY-�Kk�)I���|���� �,W�{�������|��+��� t��bNb�r1�k"����Q� i���`ĸ!�\к[�ikkN�.�}:���	<(C&{��*,;�k<.E�eѰ����n������Ն�QM�k���<`7+Xx\�A.�ң�����ź�G.�O�C�k�2b�����e������rQ�g����H��'��?�w�X�Xܹ��S��={�������tӔ)'�=p����`b��r�ȿ��׻����K�$냛�Fm��������~��]1�����������ѧ.��)>�(����0)���[����! A�P���(�PD��vuUQL��Ȃ *�"��bX̬b�,�.���,���ӹ�������g(����/��@?�<=]]u��{�p��Mx��k�.n�p�]*�wF;��H<?�ʉ�.�C��N�Y�J�>���?��N�]ش�B�g� 0�x�D�����iӦ�ZYY���6[���57n������͛7�D"ݓ�d)�r�<�Lq���M?Zl����g���NV/�����rlF�P�	8 � � ��q=7xl�� Y����q-�k!@{���,tL�����0��L(�J����c8m�H3,��a{ j��6h��X��(p��R� x�IN�\�_jN��@&�jG���Jp��3X�%�e �!��i��5��@i-�=�O\Ƕ1Fh�4G��X֤�����WF,P�UU�T�;��5�H�?ͼv@���1�/������G!Kh�5�׉��N�##*�]��0��x0g�#�K�Z5�
0M>|Ǯ
�$r��s
������?M������'�Mn&�_��<9]�H]]��p8��QG���.�أG�T.��-[��ǌ}E}}�M�L�-ytC�9A�_�v���+�pw��{2��b<{R��:�[k�z�z����-53�F'2���
��_�Ƞ@H:#�G#"��8���O��I��b<�ӦN�����VM����Y��m�R��A���g���k��F��Z�k��Ձ~����/����M��t�ر�ԩS=w�y�x��円�!�K4/b�!���gljܨ�;6H���=c�1��C� �U�i	@; �W����y۱�C8��,�J���} 	���pI�C[�0	l�����'�c&y��gF�@S;�_�٨�?4��e�; 2��l��jX�O��v��)<Ѵ��;l�x���1`� �@;Ǽ��9��JW�c���3� E��sʤ6��n}Rk�� ��/cJ&�r�!��O���3B0�0�ya[�?�R�;<�w����o�-�W�5_�t����O�c� J�FE�D[��@���Ar -��)������9$��� ��a�h!#���Z��qI"�_x���^:��%����B��ߎ=v��W\q��\nU0������yZ:������~��KKJ��;���g�}��(K��1�Զu@�Ĭ~ta���sI����֪�n>�KV"�{��>u�w:�Ͷ�>�˦�9n�e3j�8�����?Z����>�&ӌ�5���&e�fm�Ν�w�}�KJJ�-u�wg����曓���U�~x�U�Vy�O���^�9 B���j�s��yQ�/�5��!����NJc��[�Y��/n��C�9�)�: /��N �y�)�+��u� ����M����Cs6��x��0Nl�L��{ h�eQ[�yn;x��F�1�Gm�R�R�=�H�Q���]���]��
��\�\�����0'���{�ө�Ղ����ŝ����X_h����8�
�e��CP$1��ޕ@��l��  2��`G����TJME(�M@ߺm���#G>^(q{��'�{ｷ)C�0�x,)י���A�����5c6C
��0x�6���y����S�E��t��u7���r%������*�˹*//���|1|��;*s�B�����������!�K��Ga����ЇG|��'���ݹG��m�@������{llIܸ�(��x"Q��SBX�p�Bׄ�ZS'bN��wx>����o���?��­X�����M�XbL&�)��u���ݤ��2��~8f̘K.�����OKk�$c��ݩT�L���	9��O�NB� ��1�����6n�͋ Ĝ��D��f p��E�8�� �� �����ׯ)G<$�?l��|�7��w����g ��	_+^��3"��O�1���<4�Iy��Ix�ɜ �L�v����i���V�_i��<�|S �`��Ҝ�9@a$�;{O��e���]�&`��AxO&�aN}
��@~�䩄B?!SR�`jZ܇9	H����!5m
L�m�[,�V�B������*:�R
 �wlUU;�!��+W��!lU�;�s�='��qye�����'����̓�H?�SP���B)�a���	s���R���z�޽�^�z�jjj2o��F<�L��ưif2q����i�������o�:ꨝ�w�/���O>ɿ���FÑ�T�s��9�/2�t�F:��G�<�]�v�����=�?-�1y<�����}�����﬩��L]Xn�p|"�2Ķư�;��D�6���{�铳�<7�tC��������$�Ԓ�|v�Py�3�B���v�m��ʔ�t/x%�ɞ�t���3���>��#r3g�n@���ӪN76`lv tESګe)�* �|��3Ls$�1k6<2��	����N6�v�jN��E-����h��A{��Ð�� $ D��G?�ؘ��&A������/��I�;��d^�Ƴ�Indi�(�7�
�����g� -&�}�K߭҈�z���R�F�Ѐ�(��^zvY�6��1��p����c��v�{٭-L�&��[��	�$[�z���,�M���
��&��&�t�@�/�ӿ���1 �)S�H0�������&��&��IZ�z���>q�0/~`5A�!�`�f&+,,L�k�.٧O�XEEEU(?o�fi���e�V���n�5�'P�5�L6���WTt�ڭ[��8 z�I'�<�?mq��-����KL�S�M�t���߹tm������u`���w�	�+**v�f�{g.��b }�'��.{��ۻ����C��.�tBd��"��ŏa��C�N�Xq�9�^���K��jr�.]���#/ef2�h$.7�$�aU�"�Ng�n��&L�bĈ{��Ȳ�`*���i���ƆvS�N_}����M���͆��ޥU*-�Q��)S9	T�_l،�������$�a���~Eޢe��=�w�m/��`�T�˪����Zh������u 5�m� ,xl�R�����xpY��� OA�fSj�j(�P3����N Ɯ�]a��	��]Ɋ�f�����{Qk�k�Ԏq�=$��
l8�q�h��|1܍����暮��i~�is����A��0d�W��1~�HPC�q^�"AR���Rq@�EIi�����k۹Ki�9昣��_.���>������s�����y�sN-'x��.>�L�p:]��p��:v���.]+�(//���������=O</�(�iZ���^���>��xR%%%�\�~���b�
�#����~�~F:����3��o0Wmە���֥�+��:~�С���?g���s[�#��sSn=ͳ�aNIZ6E��N�qQ+�.I�S�MK4d2�������K�yD0 'a�������w��==�)U��6��R�eY[9��'M����ζ��z�7�J�2M}���9tٲe���[�*L㩴�^� �Miw
H�rSi���  (` � �a�;˪g�0��a#�z�h�wj�/ �F� 34�l��l�1���B��-&�Pk�f̼�`l�x�:��8}�&L@ǦOR�x�y�t�З�6���i>�yܮ�s�)XЕAआMP�k��N�˩�����צ��y0N��yDx@�V���> I��	��`�6���v
@��2L�`�0��C���Sψ[Tt�*�=�q���2� �!�,������/ȼ���2ˑ�As9�,v;�ܛd���G@�yѮ]j;t��c��m���n׮lCyy�*�++0�DiϞ �_�\��n/��b�{�7;�H�i�F��|(�0�@�#mJ��^z�o�v�TY���w���f�� :����/w]���JS��R��%���f�EQA���D��-U�"�pf_���'�tC��/�Y��{��������n��K�YmHn�Ys��p8�?~��s�=wo��C�T��L&s~,�8i�$��_JM(mT�k]7k���( F�4��`�$�b���.L�،�=������'�͸@�Z�g�P ���aZ���:�a͙>�)�!�'�	������wZ)�>6u���;�C��]�\��re�T>un�4)Ss���h��X)0�g���\�{q^���4|��)d�\�y����88�5`�Eih*�
����mR��� F��BA�Im�-�5�. ���6��c�; ��8�����u�,|n���m[`
?��I��2���!lӦMor��B��]�GL!��c�;�
��P^(\RVZ۾]��]�~YQ�eU��6[��EE�T0Xݓ�v(p����R�~n�J6��"�㹀�Թs�=��uٸq�P�\U���-3Т �ڲſ���N��l������D��hX��n��x��9Du8*�(ah[|ݺ��MWߧ�����M�|3fL�e�晁@�36�XT��/���Qhz���اO��w�y�#{�=kR��E�B��^{�5'�tI��f����%66X6�yRC����fn&U�g�#|� c���?5a�2�6�$��Z��dc#[c`�ۦ/ �c�?}� ;00�	R 0L}
;M�p�[��_j�$�Q��K6�nvM��L0�O�s��9
�b�{\GM�&|��o6l�&}�/��S�"���O͘&h|��an~��Ν���A��� �	C�0^��%߀��|HD���`��W^�^>�[ar(č7�(�@�/Y��:9Nxv���PBj��]�!�P��t&J����;w��m�x�[�.�())�q�Bq��i	��݁$�֭M�<y���[oH��m>�u�8�~�ڷɔ�)[z�Y��p�1�l����F��ѭUO/��;�[nj'�Ө�X�~/��BNI�D$����w��:g\�Gm�բ.^�PŒ�-��ɘ�:�T��a��O �ծV�����좋.ʙo?W���mײ��p��V��qA,k3k�,�2��d�O��J�w�"�)�w~�*PB_'	Q -IB2M�a��I".soO��*iv!�N��&G;>c��n���)�~$'����@H൬�F-��� ~�~�� N�Z7��4��KA�k`׼q^�r�\�c�� �S����KKڥ��y��Ln�y���}�d�S�f��'�$�s��8_�&@SHPV��.۴�����&��ՁadJ`T�u(�P�g�e�AO����?�SN9E�Cw{Tdƺu��̻���3�2�	������r�����Ҳ6��۷�Xڦ��?��JJJ���獴k��'������u�-��Ē��R��(݊u���D;��;v괣{�n�_|�m�.w?N�[ӹ-JC���X�&��.
6D�$��H��	��)|ȓ,4��x�a�g���猳n��)��\��ͯիW��?gxmu�,���:�0����vfY֎:,�����ݛ��x<|d2������P�ٳg���A�+⊕OWU���}��P����    IDAT��`֬Y#�?d��bΡ�c�f2���ua�5��eBl2 ���"I��e�"tL �@��}p��&JBI}�^q/h��;�먉����T�ƹݔNM����ϡ]�%��ߙ���A�r��0�4��-�~R�G����ǽp-��07�1'��B۠� �п�q3A�_g��`��cE�h�B����fv
 �������0�@D"Қ�� f���7O�E�xN0W?�x���a�2��у�`��0iۮm]ǎ�ҥ��ڶ��
}��z�P(VYY�2ϴ◵�r_<��߬[��m(� ��ˋ�k^H�`h۶��;nԨ���R��xz��Z���/^|��V�W��.�-YS#���dO  �OiST�z�.��z�Ӈ�����r�^�dqŢE�߭���ǃ�GX��B(�rN�=����?�⫮�j�-���� !�gn�tj3M�<�0�0޿X�Ҥ#q��XT$ݰ�Z�J�@'[��O�C���¯�gϞD�i"�5�ɜ�o�5Dh�X3��	�,�{�`���#���� Fa �=~��ɮG�̂�1� �$KsO@���~� o7�3T
בOw}Ԍ>������(L�L���8,|漐؇��5sZ"�&�<���
�d�X��lz	X7�	����9����E
�Z�y�e�DL�=��\��P�������@;������
�HKp������QqM��k�֥sEm��X߹K���������Ք���B�P�G��?�7�K���SO�/���y�d�]�r,�+��᫰��>,������3gU3ɱ��{�H@G�W/�"?����̔j��La"�(T�_ܐU�|�͞n�g��Ǌ���a�n;�jG��4+��җ�le��B��@ ��m��v[߾}�Zڂ�?�e9���3�^�]�X������]3�P�;��rSdb��~�GW�e6i���2Q�a�4*��ڵk�QG�d&G[8�`^u\���n�e�eX���8��}�9@�q� mlRB <Ԫ�sKP8h�5j�C�Qs%i�. ��~�es�O�!�Q#�=x,���ZE�M5�!�п�\�� �$'$,�_��c�&� }"��̺�h2���G�h)�z���1?8k�5�=�����t%p��a�����' �M�Rn�~������TB��s#����e9��w����Bu�|wm߾�ӄ�s�������?x�~��{ �ϯ�疿'���B�׽�4��&~�i��%��ڭ3�"#\�`A��������8� �O�F�I���F�Ң�V����_}��s�/Y�h�G}|��1��d2>�ء���	�d�N��9�3.��曑s~�`q666�p��ݞ�y.Z��x�駥��ￗ �d�-���az��q��.��$�Q0����=�h�_�g�h�� �@{��QC�1 66ml��t�N�9d��@����D6Ip;�Em�4�ʍ��mJƂ�2�̹�7��9n������إ�(�"h���C˥pa����8��.��1I
ǌ�Ÿ9�X'�G�� �η���>�}����S���&���[B+�qo�g�K�<X3�N�v��&��Na��L���z�8�����%�:��P>��H%S����������9�ݭ��/�؇~�f�����j��x<�����)k\Ui������¥]t������Z���[�-Z,�K-��E��W���u"�dC�<B�"�6D]<%�n�NWE���c.�_t�������ߟ����8�n8&�=�tJ0�/???�t:_�8q�MC��֢����9˲��������UWW�#al�m�^n��ĕ��� �N�RH,C��Z/5Nf��&��� r��t\-�Lc�����R;��P���IȂ��M�v�'� Ɋ~c 
��ش�=ڷ��E{l��jj�v�.5o���#��(��d5��97��q
 �Ti��@�w�K�]s��Z�/�J�2��Ve��}T$�e}�r<<pֆ���SF)`�9�@B�
և�<�9����?r�c �cz*-\!R��8�4�����Ksq6�i�?�#�9B��o�^�����30y����y�-��#	��
�ĳ�8����t��q�5�\��>2\�����;x�'�x����/�ɆF)��`���aN����X�n�{��t�a��\M�K/-������t9G꺞'�Xh��M��Tы�����1u�Խ�N�c�	�a��y���e��{���~�L�dg�Lr��O`�9���H�R*��4����t�x�H��Pb�:�%�.�f�W����,ւ��.���O!��8���T��3I;��N�F�M6�y9�ym�8}�6�h6f���u�4h��}���m`���nZQ��w��s�vi�ǽ)8�g��c���
�* {Zh����Vh�ۅ>��$>{ ��9�H�1L�[|��:����Jj��C��;T�C�Ý�M�5=��Ҷm�/s����^��t�S��X[w�)���j*Ҁ�d���������7�>��.�(w�=��9��}nр^��䭧���_S7�L�K��/��%��L��dJTg̝���2���憎:*g��믿��Ͼ�l���>�N:�r;3)`�H$�v�Q�F_y�{E�eE�E��i~��w�h��p���⣏>� �m(���ƪ�c�Tύ���a &'A����ZӤIO��V�R�[����1�X#�M-B�/Ʈ�i֧��)����Kp'��1�+M�9��?^C�%���욹�׎�O��i��wuZhݠ���+�?���Nf:-,'�05��l��V����
�a~�צ� �2�*��6I��=ޏ���g ߣM\�pF��6A�x�⢋.p��T�U)t�����Ec3�p?�''}�����f̘��W��K2��2R�7�;��9G�P���{ş~w�e�铻����f�tL��������AH��N$E�P���.�iC�RiQ�J�X(������)7!��d��_˗//�7��X�r��U
@�&��`c��-M�ꊊ�_s�5w:��W�,�aƐD"�PsX �M�� \`��F��� ���H$Tf4jsd.c�&N`õv-�[�* fX <@���
Oc�m
]Lˌr4�b��1���Ih  }(H���B
ӤR������f�`<ԤI|��۩5s>0O��N��Na�`N@����}�V�xO�}fMq�0v�Cm�*v�XJ��~���oZ�7��!a<Xkj�vR��s��P8��@�
���n�O���r�'Z~�g���#G�)<H�
�X"!Ae]�3��WŢ���t�b7o%{ts��y�i�nj�i�4���"�ƒ*U/ ���y���;i�o{��{����ηx@�^�2���ţK����V��%D2h�^��2����"iZb��ׇ��=�w���i�����N���?�x�if�84��	Bذq0	�.�k�a�v��w߽\�4�j���D�LF��pjg%�I'��-Y�D<��hQ�
�|� P�妖�M�&r!Ρٙ>h�R��&�� Su��Ijӌ'��`/ʂLn���ǵb�v,���~F�v������%����Q�$�>\*���L����Ӕ��	(���PY1�4��8��h��;��|�m7G����@���дM`&c�q_�cG8_vaB���ETp����3g�z�/��V&��l��0���Ը�;�}��m���['p�_��?�r��R���(�"��y�H4�`:�پ}�}�s۾5k֬>�,[�`*e.̌��MZD\��+�4??�� ?��+�^=����m�[_�Z�t��O?��G�=7�{^��R�9����X"c���<�n�K���\[�������֩SS��9۫W�̞sǹ��S��������Tnv�2��^\no�!+�����F�0����ҖeY�h4z��I�r:���x����{��s�\R�t���
&xl���	���$Ɏ���灌�kP��0&�0=�\�lni��t�����6&�!�m�z���O�u	�4���N;��1�� �~��'eV�E��g�?k�01
v ����w�=�% ��MM��3�����:ƋS ��L��dD�G�b �3�.���v�b� ���y�<G���
M<a*��n*�%��#�����_c�A�ft=��7f�hѷ�R~�������vWMu��i#sk��]��'���v�ƍn��֛6m�����*��J&�P��(,̗���y?=rР�7^{��6-q<{��������<u������)�C(��XBhȦ�u	��;����~�:bB.S�>��_:=��#t9]���|��'����b�1$�F^_߈�{g�n]w��s�8�VozO$������L�pb�ݼy��ӟ�$vlWY��v�C��ܥ}�JrBs+Id� ���s��H�LU ^�} ����#[�On��~�)ډn��g� �`�y�`���q�o/��Jk�R�]3Ù=���@l�Ԉ9G$~Q��)ܾ���Ŕ	T�]�sK��4�+��" b�${�9F&��;�؅�k��9w$��I���~ r�q_�s����q�c��t��i%4���u��၆b�G�i�G7�L�7�1l�)A�!��bASS�=G����)�;pgyy�-q����4���%�,y��d�`��1F�!��NCY�6�f�Es�;�8EN������������}����,��E��q��B3��҄��62"ei�&��.�V�c�{O?��\���7��o��f^0/x6;��9U�/�Zߪx������tЭ��x�N9���I��[��FNM�Rw�n��f�7�xC���r>"a�����=���#I���	�k� r>#� M����d�Ӭ�ID�5�q=��f��P�V�rIS3@}�ྸM�L@C�19r�菧�A���_K߲�W�s�v9��	����;@k 6a��� h��4}�h.&}�o�`l��SP`Ȗg8�'���>�}�y��c�f�1��K(!��g�v �ƨuQu��>p�]�����+���^'j(@���lu�T:�Y"���S�+������T�9���o��u��!�2as�=*����c3v���/��/��{�[�W�_z�����lc9��DJ��n��+��No@l�Q-Ҿ��i��w;~��&ݘ3"��\4w��E���L�l��#�����<�ab������?qƈ��Ǐ��Y�_�.�X�<����q{/�,�@����c���_~Y$�PE�;��=���e1���N�"��\���������@A�k��yl�*k�_nBv �M�`�kJXgl` !����w;��ٜ �~�Z�Ӯ�7���	�4��3�i�
A4�Sg��1��;���/�%@����8�e2j�' 
x����D|���?�5�\�Fp�g'�Q��s��L�d:�ɀ�q9�R�B��v*"�k׮��/R_1v�w�4������@jiS8Q���J$Sy<b~^^�}��mY�`A�g����T*uh2��fr�p�����5M{�����8����v����{�cY~�����듷$�sKLG�/�#U鼐�ݦS��R"�q���,<��s�1"gf�t]������#�ɔ�;I�q)�06$l� ���XXT�ܘ�c��tR�ϖ��2t}^(�K �����͓uӥ)6���E����
p�;��v�,f��1������W �X 43O;�
�� \��f&8����t��=e�P���H63\Ks2Ǆ1����5i|�s��-���4g@)P�g�`N��] ���ڦ����7$��*B�VN`�Z0Y�ѐ��%FI�㶛�M���`��}�y�sCA��T�W�A��!�%�0l�� $�y~q���7弧��Wk��-�Z�L�&�iS�����hW�ZU2���FÑ�k��p��L02 s�5��YY���)Sn�W��|��(@Ǽ��9󈍫>�s�P� W4&�dLx���l9D��@�44��e�*g�3we�;�=o������,��F��t�ƍ�A�7��A�p9�"�R ����~]:�;aE���u��Z�ⷲ�pi<j�u�\��`$�i?�`�Y�<�+R���`���a�~iv%��Ԍ�8�̘k�*6�`���vc2�����V�͟� �&yƂӷMR ��h6�yrS�j�Ԭ	�v�'�`eg�S�i.P+�?�g�;M�s{Ԥ)��O���Vd2���8���G[4{3m��I	bph�5 h��0�����s�З��B(�SS�Rn��ڰ��7����/{�����r��1��]�[LC��ttjտϟ�!L�6��믽��������L �����`8?��o/��]'�|�����~��� =�jy�k����N]��L���i��j�y��pd�ˈH<-�.G�ʙY�����z�؜���x�6�7�*�0Ƙ�Ym��?}ހ�7�D$8x��5�>v��ɓ��='�����o�$��nl��۶M��
Гr��y�t�R��J���v�����v-}٬=NM�0��T�zk�z���K�M��1��zQcg�U���������q?��f<� D���*L*Ԕǝ�.��B �A�� ��L�e���y �'A��j�0�����R�b�
4��-��S��R�������;���Z*�k�fO�z�"&��Bյ�,3����*�R�;mXS��d�K�$���*�g��p��ø����p��7r��>m��x<1*�N�9����.��Ѯl����8�+'N���˿�G��S�8@��W?�h���^�U��o�.�&�.a��u��C8��\bGc�����S����t��ۺ;'�����ӻ��ފ�5M�N�}��z��"+�E"�x۶m�:��o��K6�O-�]˲�X�lCO���x:��C�^\֔E�+LJ����ӗ�yd
Of/�a3 H�H���L2�u�v���]��qo~a�(�����]j�d���vS<�u�r�lv w;�Aȃo��y����Y����<nHZ/h>���@˴��f'��d�l����8jϴ2�Mf����k������P6
�?�+hw8�@��������|���f�$>�"���
���d�w����W�q��,�d8��4WS� !ĺ�"�OϏ%_����-���R�0uҤ��~�ra:�>k��J+�k��KAAA8//oј�����l��Wo�tk���9#�e��)�kHhB$�­)����NQ�I$��x�;�w~��+/�_��ԃ_x�	��5�Ģ�J<����UR\�T�"�V�iS�ܕW]u{k'�TUUuw���~�x<�RZ"|�ub�_|�E�b�P�x�i��p5�*0�v�;	_�ہ  0�R�Fr0��<@��Hb�<����hFs?�KS-}�4���N�h���Sh!`�5�c�	���Mm��(���!bL�B!��NP�;�k'��<��y|Ͼ�5��-����.
{(����r�)k��YO�k}�� ��5�~�/-6nE`Df2	�Y��������F��dbw{US2Q�u]�K%S�����������ٰhŊ�f�}�]55��4Y@�O
D*KVQa�g��5~��;?���l��H@ǲmY���[[:�4a�]&!W2-DZ��UG6yH�0E4)�ר��>�z����sB�ꫯ���ᅗo۾�*���<� �����$�@`c���Ϟ0a�Sݺuk�%-��46�J�����aC�D�(�}���w��l������,3�Z3A�aY4�Z<#{"�
94e��Ž�t�"5Jh�_�9���&�Fm7'�Hڲ�}�|�w?��$l1T��d�7��$�;��)�Ph���$�q�Dh׾��qC��v����E���s���9�+I�L�C�}d��_ :-)�E�����/�8h�:��c�jǼ ����t�G��}    IDAT�FZ8P�y�d��l��#�\�!��J��7�Xef2�KJھ���`?���2e�з�x��n��'�����T�W�*��`]~��˯;w�v�sfy����:�`�=�Y��?��hX�IN�@��rZB��"��.Bu�Y�hW�ҁ'�r[���ݼ���-͟?��3�<=��ε,� �[ŞuIj^0_j�a��C�N��o~�����զ���b��j��/��4� U�(�;{ٲeҧ0E�=h�4�K-
�M�40��Xj�43���,Ik��b�	B�
l� � �v����.�6��i	`A��L􁓡N_7� �(�1F��9�k� ǹa���y�]�ߓ������}�?]��eXf֍r�s�7�c:�	� �y
HX7��$��]B+�=����x�<���J!����o~3JV�S���N���� ��X��� 5n�3c������ߗ�Զ�=���]\������G��~#i��� S{����?�?���&M�,W��v��أ�q���7<p�kgÕ����/����uk�pdD��AH$tC�S���7�mK�=��jr�pL�8�r�'+ge2��N��MS�d���C<����D�I������׎3�Uǧ74TH'�Yn�k06�T*)"1U�	��O?�T�!���H��Sk$�wl7�- @� 
�b�8���m�6��� ,���	h�P��̰,��ч�������ڷly=���O`$��fh��i�oJF35���ϩ�qo�ߜ�(���4s��C[ �������1�kȸry-"R�Β�(�0�@nD�B�� �p
�+R����q�9g�nݺ5�qo�$Q�A�$�g�����H��yM��]V���\�	{b���ա?���+׮�z�eY� ���E�������,+-�?����ýuO��_��{4�c��.Y���7ߝ�n8��˓�K&��L]3�������hZ�'RV"����Y'���5��"���^�z�{�왧l۱}�i�)A��pF��T��D*�h,))yq���SO?��M��SKh��ڪ��Nm����_�%M�ԑ���?%���?��n�J/M���Η�>UV7(� &{��'H��F_/�������!D`]��Ì�p-2�q˨�ٱHl��A��$`��?	�B��u��@6��1�iZ��Щ��z�G�>}�M2�q��:��ǎ�}`��DY���}�&ϒ��0��B�����gt�,|Zgh5 ��3��Lp2�!��%.��bѵK�l:aU��fv�x�|� �B�4�����VZ���}����?��AO=�$�p����ZS�ę>?2�Eqq�����:��c&\w�����fo���X���t��m���]fXG� �s<����˩	-��[�6Ƅ�o�>���FL>x��ks��˞|��'�����:���l\�1e4���26���;�	ysڵk�d�ر����Jq���.L1:c��5M+N�*�: yÆb�2�4uV��F��l$Y�^ �)T-���瑸F "��Ә!=7|$���m����p?��	�La�n�&����kN��/�Xvr���0B %`��P.	������NM�`,<��0B ��e�v"h�z��qn���0�Rh�L�����G��?�����h ���8{8�
��1Ы���e���^x��d@8U�EU��5j�0�u[_����W�\QQQÿ���}��g�w�q��?n?۲�R{�W���2����6��is�u���ɾ}�����i�cl������~pFx�)e�t���2�éԺ����P���R"&\��2v%%���z´��Y(۟���N+�~sb}C��.��Hjc�b_y��)_z�l�]Ϟ=���k�ښ�Τ��>�dl�%�a�ӕL"y�$'���~[�[E�\�Z%7�ɕ&x������M���F�1�/̷��|�������$�ײ�U��!T�/��0�	�c ��i!`f;%�(=S���M�?��+�P�1|��Px� @5�i'�5���LH� #��N ���Y�/��'��o`(�4��Ϝ��Ԝ@�I��IKN��=�Y�DY��!|��PC</��z��%����?�p���رc�������o��,�=mڴӖ/_~��=�|)akEb�
�b���a�N�t��W�Z�➲���1��^|�����ZM����U����HŅ��T��ސ�Ӗ�&tw8E,��hth��	�����3g��k���뿙�J�'#�96#�qg4	��e�
4ClD�H��~��M?~������=�A�9�D�X���x,9��u�qCӥiy�ʕ�_��A"���Ti~�X�0Iiz&�!�������L� f���4O�\f��anX/�$66܃���`?;�Q�&��M�������LG�����ڵxj��?CԨ}S������k3Y3�:��f~�}���9xG[��j*RC�	Io�'��NX���V�������iq�p��x�ǧJ�~ġ�������G�9�h�*W�J~���D0�����^�L'��ѣ����������̙3�ԍ!�d���
���)��?���'^~����J'�{�j3�j 3����n[��΢drH��b��t��٣��Ws	�p��#Y�L��pu��Y�y�k�rh*:�3O����af��ij؜�HT�����$��z�p�]?�c&^x�U����K������D	��$3*���W^yE�*A~n�@h2Ӻ�GXY�@� ȍ�&a���4]���ۥ�E9M�1�� �d(�
k$p�@_4���=h֦��'I~v�}Gh�|�{�o�$�4s�A�w{.z9�
��ځc談is���s���{c��G@���qI{��O9���V����Ζ��5�v�@��Gu�6�d��yd ���p�d���1��7������#�zE�I׾���~���;��n݆1�xb?h��*�%�M@>Ĝ������x��+�9r��-�!jU�nm��{f��Ab󏳋�zo�,l��0#\�&�<~�΀Vn�p&#j2F,V��|��M?���i̐��歷�*��=g�~suuU�.��y}Ai_r:���k��h��L��\����a���"�He]]�L��{,�h��SM5�ʶ|�[R�c�N�r3�g^P�S���EM��d�����<�8j�J`P�2�=�@Լ�?4��]#���"��d8�ڙ��Ǘ=|�}�fJ�� K�m0�� ��?烦j
.�`�\
�#�����?��k��GR����c��>�H!��bG?��rKSdQ��H'j�M�{�G��	vqAa���SOGy��<d,ţ���r��z�'�
�e9OQUU���U�<p���;w���m+�`�����v�|#m�F]H�5�����<ʕ�7=^��>��3�^�ʧe�^�t����W������[v�i�rwr S6g##|�Z!�.�q;����H���3%�o�|��]�ŧ?��Cm-z�R+c^��۫е�p��Rˡƞ1,��%�EE��<t��7]���D����W�y���e���cq�"��J\ ��^zI c%H�T9Z�G���;��w[iQj�j�:h��3N� ��4G�v�Z�������E�J��дO�%Q�&f� ?3D�>d�T)`48H��sH���%���1Ѫ�1�|��AK�0�-�9����'��1�$��%���54�"�A�����Km<Ƈ4����Jm&�~���9��U�}&�irke3I�t�L}?���k�w���A���(��V������}[493���y���Jͦd�y ���]z��p�	�6)����Zĩ��1�k�<���%������fa��-R��p ���-��pz=�>��/3�&����C�8}N�s��a>����[���7Dc����d�`�-���ƭj4��#�Ͳ�z����Yg�9yܸq�2Ĳ��͛7���@φ�Z��XVSS-�x�	��\�ư��M$�a*  ��5m���m�<��`QY����Hm�Z�� UU2_4�@��,���fHB�' ډm�s%;�̨�77��	����@���v�-$����;$�!���x
I���q|���m8�c��r̖"�Z���������f~cB�n]*�駟.���+��0u)�b��Ú�$�i����O��,����_�"v��	�Z��ƇO����L��=�tZZL0����P��M�@v��%��:�'N^߂���w�U:V��?���ݏ�h���n��-c
o���"��D:e
�p�DF����S���>��I'U���������ޟ�_5fN�4-/m(�46BH� �a�j�UQ4S�xܞ�]4j�^�*<�e��V]G�))))�|�c�26�Y��_�*6n�(?+�Q�MM$�M�ƨ]�p.5o�5A^�4!u�K�1�#� ,�g[
"�g��e3 L�h�!�I��/��OY���@�Fl�%���}�k
4v���1��7�4Y��Μ�f-�Ǭ%�>w��mMLw�m�
@F<�yZ2B�ˑ�m+w���=n�sG�z�>H�~�i���>_��B4����G;�������1bĊ\����v|���W^y�ު�;�N�i��WR)9�ҍ�'�廊�}��;��q���֣G�}���Б�x�	�D���Om2ڀ�i	�%d(��1��_-OdR�9}"�J;M����=0`İ�
�Y-�1c.=�����nƐh<�((�T@� ��2,�'n�#γZs���8c�ԫ��*�Y544t۸qÍB�s+**��t�)�7���>O>��d��a��d�l=u;�̮�RC��� ���� ��wvm�!b�ğ-I �I����NM�!���Uܴʶ�?��ĸ/|��5u���6�R��D'1Z2��$�Qر�H\�D��%@�	��1��h} ��{�O��P[P����_Y#q��z�^=řg�)���QZE�]�ˉ��j����Zq <zm]݇��5�<�MM��1����ի�Ϛ5kZMM������2n_W�D.��R._����y�9rd�B~[F�Q]i���UX�reh�3Ϟfl�<��tv/�2"��
͑��y���p	���Bw�S�PpUA����`��Z��\�&2��w߽��a��d:yX(�j�k�G�pYq�L���L`B��/�_~�i�N3fL�,�Z__�����{��v��> �rt, B��X��	�i�@�Qd*j���rc'x�������Ȩ��5��&}j�(P�'����dM�Ibȡ`�
 �7�&�s����)l0����t�5v��X|gO����8���	���U
=@i^ǵ��o����!O��J�#I��Qy���N��.���^�I\I�����M��tZO��a��{�u��Ͳ��H.~�{r�!�4i҈������[���`��;�4e�v�޼�T4�L擁�n������n�}oՀ�E[�ti�ϟqLQ}슲�(w��"��i��f	�/ ҉�8�"e
Q�2b����e�|�a����M�_|1��c=y���aUiU?"�/ۧ
`������UU����ŗ^|��Q�Z���s��#W����+{�����E�p����x��<!�>t�4@��n?;�ZinL�ls
4��c���*bh6Y�=
4��5[��	�h�&jj�c&�#e~Vn��ߡ�	�d�s< ?��*�ܥ�R�l�o�������(�����!�2I�E[t%����e�[f���J���oX�s�):� ��zq��cA���yf{�p�������p:V%b���mU����{:0,Y���E�ͫ��:��v�Ҩ��T�YK3�%�4�"?�;v�9�`��s�k���:&�Ç�w���On	�6����+�D#e�3NK8�.��^��.�)��0#�¼���;w�g��u괫��n\��K��,^��Ⱥ��	FZ�!���.�6-�,M�D4�$9�H��΀�������	W�ۍ�iMY��ںu�Q�X��@�`0���u{��iK��o˗/���&$�]	?��8��@鳥i�D)�8HY���M�J�B�;h�4o��e����/�k����j�v-� E��9�h�V ��wi�J@��f����p�l�\ ����v
$�-$���
;��R���OF	����laQ���SĈ�{�������ay����4��K�JW��-�$���4��
}XRR�K[�����X�vm��n�mJUUՙ�D��\w]i�(C�g�q���P$�q�ɧ�|�e���?��Ks8{�c�^�<�2��_3����EN��Lą����W�]�-�05E��m���t8��ɽ��^��(ғO>���G�0��_][W��%K�P(��/�g�$�X4Vݶ��s���_��|�9|��צ-����W0}�n'h�����R�� ��\�Y�Fn��(����*�_�,����&Rە��Jm�*T�.5[}�s{; x_j��A��KS4�j���M`���6W��k�v���6��h��6M-��͔�v^���OK��=��{Q�@�H��YM�A�a���J1h� ѹs'�G���;+�:H�@��}��Sakh���̌��Եۃ�������B���_BFgΜy�;�3�����S��>,�4p(��	C�/{��1cƽ���k���}�@�V�p=��3��5��=��Ê5�ӕL	���i8a�,�A�.M��)��r4&��Z1��^��u��ƴh��|�h�0.KDc��l�ΐ�`0$5��ƈ�'���Z������L�0a�׭-�6�D"|H4����`+��e���j�B.����X��GҊQUU%7t��<E�SU��~u�	[j�UG��J� �>[�ϋ�TM �:A��L�&�Rc'!���ݬ�c��P��~�l�8C��&-���C�m��5f��{c\�磯0�ة��/�v�`���-�F��eY��s���}���{��%�~�᢬�H��5�vO�M��v��.}� �۝�'������ҷ���� �>�l��{������dҗ�(P���5U�������G/�����x�?�߰��_k�@�W�\z}��A������vo")4���Bs���҄���n���.j}��pA�{]�s�!}��ɕ��B.�>���!����t�-�����J�J{��&�eY�^�����O��⋿*//ߕv��z�v�}��'���XtB4�8.��Ya~ �ŋ�am ��� �s`��ixUz/	�������n��0��}��Ӝno�EN��9����k�v�-Ծ�6�p��^8Nm�KB-�n��f�僧�?d�SӖ	F�Y���L�}���<�.�H?y0(�0ӲҸz��xFWE@�]���5�L�$9P(2B$e	��X��|탢��}�����"L�w�u�-[�n='�L�S�f6������^3�{��\3v�5_�Ɵ���r0{�c����z���<u��������E[ӓ��9e�ff���Ad�����-�H]��������{��"W�>���o��浱D�7²�2�,8����K�����t�b�x|����袋Vr�!�j#CA]�+c��UUUU��*`Q	H��n���_�"�m�&5��a�W�W��Ԑ	J���NKB�����<���wH�05H (���3!�V;1��:�ή���D��h��q?���:2֩Sx��盃-�_�3懂	�dp��{
v����sHaﰪ��d"&:���%�����7%b%<�W�i�5���T~�D}C��D"�@��6/�K��?#E��~�k���']�{"�s��>2������m(/�}YY����Mx,��.r�m{e�{�c��z�ɶ�>�꥾��妶�EA��H&.ܚ�<izO�enfD���`�k��~G6���C��*+U��n~�_~��k�����d����Y��S�Č����4�L�{�4ͯ;�9�\r�[}���Yb��<��9˲��t�GCC��d2J9�@    IDATy���@�I�r8e�:��"U,��?�ݏL`b�u���E����O0o��&[��n'�Q�'�+sӜ ��q_�Y� ��m����Ԗ	�jx��3�	��� �����O�����:�'-$�1r �J�]�)��$�Ő 0�<;]ٲ����#�ӆQ�FV�������**�i��ۏjɒ%=/^<'���<j�`r����Z@�7�a�����}�I����4꿵[��'핀�)�`���6��r����w��U�6�"껥�,U0�!t�JZ"c9���:�ll(�[^1��i;`]�@}�ܹ���ҋ��>����=��X\i�%�M5��_�oP^���������E�w�'�tҖ_����w�,�b��m'&��+
K��xZe�A�w��E<46'|O2�݄n��uS�z��L�NB�;hRs���}� 2��&g�C`���\C�9�+}���l�7�������D;�I���Q ����fz�����>�|F��-ѵ��##��v�ڈ3��.��,㞒��jk����Ϲ�~���ތ���o�qU�6mZe����KZ�~}�w�q˷�~;��v����+'�&׭�N�ǝ���_կߡ��<y�*\��ƶ�5{-�c�oϛ�m��_S�1Gy�ɲ<3#<�)�T��#�TZzC�ґ+�)�.��r:���͊A�r�_j���r�0-�;w�%�=s�д��D�0UU,��Õ�+C�r����E-��N�7u�����#G�9��s[]x�eY�pݑ۶�!??��C��_�z�j���t��=#5u���Nɴ�T1�6�'�!X��-�3���p&�/��`fx�Ń��)��O��ݤ��YB�O���b&v�G�)X�Ԇ6a���̱S��g� �����*�G\g�wn08j� o��BG�=��ӆ��i���9&Гs;}�vAP���/���\�1�X��ڠi����aki�3�O�>��޻/�JU��AѮwM�~�~϶�?ϸ�;w*�� �Հ�5zm�̞?�Y;�_�ǋ�C��"���<�W���|�J���Hx|��!�VIѧ��]f>��On������ʛ�^i�\�ҍ��TR8�4��
Y� .����HHpJ�RU�ڵ}�أ��y�9�|SQQ��C�����ey��i�<I�ӝ��4	����;�H�E$�dR�;M�����i��P��a��eٓ��ݤ�Mh٤-0�Km�@���g �Ԛ�n�p���͌)P���Q.hL2iK��(��vS�a*���a䵷k�v��E{����Ob53���mQh Ü�P8�����`�S{�I��ە�GU���q���ݻwC��B�X��n��_����=O��t|c��_�n.�ԳgΊ)�[�r��/��u���sOp8�P�<G�{��d��Z,?T��Q�O9r�w{��uso����6kV�M�����5�(�X���0O���u9E��n�ڱ�tI�{��Hke%ϔ�?|�Y����I9�G�s��K��(����@���%pC�aYK��R�.C�� K@��D���ͧ�+�}�e��>��TR�V��k;UU՝���K=sP^^����'���_~ElݺUd� �sg��e�PT݃Vh�M���ӻ��J-�4~����'�1c	g�1r�b�+`�o_�k�ČԦ���H�����,�u����1i&73�)�P�����$�9Tv4u��}h�v��v׃�"|ف�n�'����{!׺<OSy�i^O�U� �/**�ւ�B)��w�9�K�.*嬩�[mC[2���5M�r�������R�ԪD<�h��tEyyyM+z�s6�-k�O�5��m۶�.��dF',Kȅ��hD��H�/[O~��G�aʔ)�*T7g�����5t��;3g����S�#��:�B�ꝢMa�0SIiZ����%4�W$S$�Q��ף�ڼ����v���ۚ��	�g?��F�[[S����J.��6T5�@^^���M~d�4�f�\��ό<�'N=��rѿ_������D"�[d27�#���(i��o����o7l���\��Uz
D e��$ g��41�]^G2���9��Ժ��;%`;� k/:"}�Z�)TN>S�,���l�&��ɗ�M��6�oY˖廩���N����������9~�v��c~�	@�n��� ��=�,e��d\j~�p�v�aÆ�C�+y���<P
V)��>IKE6g����f��[�T��6m�������������B!De2��3(�QF>s�)�ȵ�����<p�����K����qK9s��Vb���}�?_;��̜2�P��Q}��
\�攚�S@���������o�%���=~Ai�.��,��o��瞻�6���d"~@*�rJ2~��t��DaB�R��|��K۔�u�)��2d��֖�	�b׬Y�3?���T"=�����C�^D,Z��X�~}S�(˘��L�b�8i�J����d�R&k��k�=�뺪��O��v�.[��&w;���ĩ@�	�`h�IS�0``��o)C(3�G7$���8q�c;�M��lٖ,Y������}�q4y�#�D���u����)��������廯}��]����I)^;��x�(�w����� O����,{q�%�q��ٶ�>��B�s��.w��G/:^���$7�Z��e{��|���<H�r��䆒�h}�5.>�'Ǆ�as�R��7o\}�U".�ID��g�V���!^,װ,�>x�䩧$�~���+PD�:��IY�zuӷ���oَ}���H=C8w^���	�C�k�P(��#ϼ��~��>8��o�$d�fD诛�5��?���;�X¥�\�D6sT$�$	d&A@QS��	�. W�~�a�T�$�n�E7_�t7k��.6�*}�G��<~�s���O$A�����+RP|٢����gw�%�d�5s��ht�������|d۔)SƝ��СC��̧��=~�kf8n@r�����D�X��H���U��us�>#\�K���"���%w��,y���DW��&�fyk�s�{�[H����x^�ˏ���{/��~�k�uA�����������~�h���·��3?n�[��Wz�ͤ�gc�^wͺ.ʞ�6��1s:��=�V���#��\*sv���1���@�� �������%%�M�xyAd������xgGǁO�R�q����ൺ�łU����A&��y�e���׿�o/Ѣ� ��fc"��e*V��嶮�;?���l�<���  0�' ��}�֘���tt\f=�
��Ϟ�9˗�=q�-[��Çf:t�s#���)�t*�.:dY�;�~a
2�f!g	���3g���뮻�[n���x+G�lޣG�6�R����}pp`��	b�W��������EB��@.��	�qk�R�o�`|\�q�Lq��o��s<��'���퓹O��z�2�c�_V:��L�^<�	����=�
8;~�>�㻯C?:Qn�-�^�}���/Go�_��8@��W�J�Е��
�0sV�p���X/R�=Z��{P��0G���٬ut$1��s�٤��{I��p����~w�����s���t�!��lJ,���F -��򖖔���c�u����E�y���u�!@����2�~�����+AyW0����,0\t@�$�B:H��/\&��Sh��&�C}ͪ�n���e+�I��}�}�m㦭�ͥ�wd��*�8|��/SLp�K�,�s+�{�1v���f�UW_��뮻����}��O��*�=��m۶�"IR��ݻ5��E:;;ٙY��/�"��gmg���(�:ku��j�r5?�-T���m��b�(�ac/?87�������?��;8f-ᶘH�'���D}������d4��N~{}��~x�w����<�u�I������`��ac#��5w�W��e�������zhjj�	�o�E&. ����uQ7\E�!�aw*�^�I$���x�	J�*�IڲeK��|��O$�>���W�||�����<���dF��׼疛?���|r�up,��w"�?2w���ÓoX������Y�1� h�2��pWz8vi�h�s0%	Ҫ	]>	���笸�;������cނ���J��V?��\ںݶ��q�|�$Z���b�0�J�ry�E��t"
�9k�n���箹�q�0�XtwwW�R��g�y���o�jhx��'&̞FB�	�'t��Io�טe���[��w��➛����0����1m��J�l$�r��p���Ȃ�D�oGԮ{����cr�X `[��J�^�T���ό����s?��6�L�Otÿ�xG���-���=�����^\�Ӹ^��!Z�N�>]X�x\�k�䂄�^ ;��c(�5E;><2����_���=M�L��|��}��w�Kk�}�u�Y��uC�WxZ�xC����������KO��~��b8��������u	%>P#��,1����ɚ�/�@ te1	,�t9$9��+����-W.Z�,��O~����+�����TMkK��A�b�/ZL@������H��_��e���~a�5���7�p����/�IsG���uv��y���۷o������ T?Q��IF(�I�K��|�/���qA�.p�5�E�3U�@��k���)�b��2��.��Kt˙^2��v]a��9��J
l���	�� I�qX.Z�X��[�X�o����o�����o���a?�O,f�^����c��|W.�V�v�G�ٗ/_.�x֢�<mv?��Pu����?~�kǾ���-�)��kn:LV����`��~�_2�컇��8�h���B
�x?�E��aEQV�u�_���k���g�=�"�71;~���}ϯ}�s��_����I*V2��(H�, ����Se0u�oisP�]�䖧&�X����Ww�����O?]�r���t9rW6g�Ͳ�R�,�^��0�o��Z�	�o1*K�*�[['����o��s0�7�9����ñd2Y�{����[��{{�{�Ec�-���ȲG��g��N$��U��-w�*�Z�<�� �4��.���5PqѐM��xnu�/�v!�2��
9�����r%q.��1K�<�թ��?V|��~n��+0�Ϗ��o�$h����#���/rt�G��!Ƅ�mfo��hj�p6��_��^��+��@����}��7T�O�|��R���$����ݕ_���Lf:
�y����/d�YQe�ԍ+�������k�w}����D�or���O�vi�ĉ��Ts�+4-��"F M�{V�*�����,jֳ�#��)�Vm��|֣-�ncc�N\�r���+/Mݱc�g�}���p=~{nN�B�3�}e.\�#������ֻ��eK�x�C���*�q�����'&mٱ���7m�|pp��w;g�^��in��$0/�1:6퓚H�☈���y} �}�d��:�	�@	º� �O�1+>/���m�H���Cʵ��"&�9�^����²#/Mt��5:Q��Jq�g���gG����w�<�w��V��w`"񲴴T��`X��K�.�ٳgz�P��x���q�ڎ�L��S��il<���6�&E�� �f�ƪ�|��ff3�:��{D�V2�0���$����<�{��{Ӧ-w�S��B�^����]~��_^�>v��:I_&��c.C�:=�����6�3���خ�Wrl�n�)�펷L|������r�qԥ.`o�����ɧ��@6e~(��N��~�+������qb�om!�糿3�h�@Ä�U׬X����N6ΤcĞ��PGGG呃K7o���'ON�d2Q�v�&"�D�d�,���>q
+��LtG�/Ƃ��Y++�c��30݀0����a4&j�A�t`�9�C���YH86X�EB�^��Gxad_��5R�ǅ�~��O��3�__��{u�f��	�_Ȍ&s�'��VlG���X�̙3�+)x�y� ��c��q\��qx$e��G����.h������ի��c�3p�0OC���SH�@�ߺ�������~�on��/tڸh B/pj�޽ڳ������������&hs��
L���Y���+� ���T�.1�ӘP��j���\�6uj��a��͟z�����wu���2�� ��ZR�4�&�x\|������#��l6�k��=z�5��t���3�v�ԩ���O��۳�#=�O_���ߒ���-��к�邘}k��}��pqۮ��νX�X(q)�S��d8�0$	��0D4ہ��c|]xP�DKK��T���ө�9�0�� ��<��
p��vΆF��}"�;���|"�9Oȸ�����'���|�]��'�tO�mmm�����P]]-�o��;�2I�fs��d�Y=>���@�X>� ���|蟓��{S�d�w��^75ד����'���5{���ާ�<aw�/��& B�@�~������M�����L�7b�-qWb�倌IAX�P�v-�TBZ\��`a�T�!%��ζǧM���+�=���[0v
XԿ�oM߽s�gҙ��ux"� ��� vU���1�������ş/+r$I>��7̙?�7�x���ǧk�����_|u�ƍ?548�,�5�D�w�#�{��_c�->Q��si�"������j�`�=���e�gLP]�z"z ��!3Ql�")³�t��o =�c�}p��i8�MA����-~��?�j7U�_���W���7��_S��1ڽO�>��!
U�`ʔVX�p�h��I����V$9%1�n������G���r���_9o������_��/?*��Ll+,���U������+?��;�r�7v��i��"��0U����m��]�9z�SZ";��)���A� C�1��;6�T0$]�'c��)�V�3 ���hdcݴ�?j�~��΄������-[��q`��sΧ(L1F���R�|C�GW<>�{�$IJʒt�������\���˗w����0c��Mk�~���S:;�����KS�ԄL&Sf���q#�y��E;5��^,ES��]������u�뀝��� ���A���C�p��
u9]@�ĉ���S#C��s
z�#�o�b1h˪h�kT@�Z瞅>��}��p���a���|�<.CF�����~B�L��}��x�L�<	f̘.�CC���ܜ���<�rw��j���+*��ee�#c:Qt�����5��x�k�800��l6�Uܧxo����<c��0�/���>��|��Ύ���-�籗�.���������%�d�DJ�@�d�D�+Z�1#:��dmP�W���$��*g�F`opbݏ�^]�x�IV[�~�C;���?^����m��;�L,u]�D"ĞWB�v��"A0`bǗ���Zݒ$h�Puu��K�.}�ꫯ>��֖�q�q�o_߰aG͞=��688p����˲k��a�c��둩��QX?��q�Nm6�j��ژ�4��)�:X���fl����F'6AYu�N�@��pbdN�iH#��-tIT�s`�0��8|�19�s���G���,֍{�`��z?��w��V9^�_���C-	�-QuM���
�9s�`ss�H4��s����X�����]}��_]�f�s���;Cf���������b�t0�ٝw�s��ŋ�������v"�1���k�_5���-�P�o
�3�l"���58����-"Q%?M���f*���ʄC[*�&?6yѲue׿�k�'�9���߾����/~l`h���4gr��*\sX~����9���B4��1�ݽ�t?��s_,=\VZ�č�^��e�-99^-v��}��ǫ�[��q��Ǐ�\
�'�z���N��ʁi[`q[tB.n�mU�p%Ѧղ]Ș9�w�	�t��P"3P� 3+4��6��P� �P,`p|��%�ᔓ�>\H9U�L�5���F�t�%��$�A:�G�t	3���^tY��gbٙ/��ן���o�˝�zl[�h��455㜯ZSVV�1k֬�����}��l߾=�����Z�C    IDAT��޾;�U�5��\,<&�)���D���,]����/�u�Z��7>mq @�>����׿nݹ�묓���N��L2�Xu,Q�$OC���pD�0�H��ѐ	0$���Ɖ�ۦ�`��.?�ư��3�<S��o~=}�޽w��,Id�Z&��GiR�v<ˬ4�����>VU ���H2霧��z���i��a��e�Ϯx�Mv��z��W�O�>Q���?��ɞ�dS�R�ty��F\	�ޞ�.�`b6�Q4���&��s�'���q�&X�4H�&\�!=�5"q�U�-�8S�`��8���Ci��v2xCٜ39��(H�^f3��D��hݷ�q�e?{Iy����k�	�/֔�������y���N���D�mܸy��i�JKK�ٟ��i"�1�By����7�9�駞���8W�"��Q���s\�����L]m��?���Ӳe�3��MB6n7#B�=�fM�޵kۺv�WY\
Wdz�@DRAw�"�u�YF���u�a3&6Y�� `���#C�ە����^��Wd��Sc1\�:��#-ϬZuS��3�s%�-���0v.D�|�/ ��cb|�� Xl/�[���<�OU�wm�p4��?�x��]���X�����z�o~��[R��¡���������
ǲJR �b>��3B�5�h��9���? �׾'w�
&��� We!�	��%�2B(/��;��s�YQ%P�0�r�FJ��H�H]K�β��ê����L>z��e�*���t�EԞ�6�S�;�?��j�g����������y(�:u���ys�JK�v&��m�\f�$�]�����veI_��4����w����+�I��{���a�zYpqgƁkV��ԝw��2uS�@v�OK�~ �[��۷lh=��֏꼡B�[�dFa�r�c�Ѹ�M+�
M�T�Zǖ�:�\�]Қ:�i�'N�e��k�7�tj���k����7w8��C��2�&drYEX���T#H)ߖ-���ə:��	��ȉ$1-�!Ɣ.Y��͜=��^{����8{�L�[>�ѣG'O,=�y$~`OG���]K2����Yg;vEδK��p(=0(kٜ�l�li��Q���4g�z@2��p�%e^� C��4l�:���j�ŲH�AX��kꟻ���?R��x���$s�ȑ��t����ȑC��"�%.:���p���c�^���Dk�f^�$I�x<�jmmM�����b���@`���������pw]]]b��c���'�>�#�~d��~���k��8�HȢD-_j��s\���F��L4���>}��f^~����.a��҉������kV-���.=��kdͲgB��TZ$����nI��E|]�`�U�����U{��GSAu}��iOM[�lS�Kh��X�f͚�'�O~l8�Xh�v��<-sY��:�
� ��0p�_�H.	L�!����<=s'�]~�{��[�x�����;�x��K��x��9�H��ں�����	�]]�y*�8!�Q�Elp��V� �7�d�/����j�"��ð���ھ��YH�h�&�u��K~�;�x�m�_t�-���,���纰ض-]9�ܗ��5nB2���0����p8<�F������������m��  $��������e��9|��������zzNߡ�r��А�%@n�=^��00v~����1ق^�"�s<�|��Ж/M���?���oYN�=4bD�n=�H�u�`#����.n�R�s�L`˨�!ng�w+��Msf}o�WneKf���%lٲE}�駛^ݲ��D2�g9ۙ���J2i��� q<q��"A��DO�E�'\�g��ݶ ;��jg�$�y��I+-[�u��7c��Sl�D^��l��>r�b�����ذ�.-��rjYڄ ֯� ���Z��o%�������M�[�������W�~�ߺ�wz=|6<_�����{���$I5�����:�,g5M3YN��@����]��쮬��YU
��ҡP(�iZ�
�W#��_�����{���q,�S�U�$�j���P0��g����_q�r�;/�9}�C#B����;׭�ٽf����w2���Y�X�q�\�� a�TA=x4I�EYQ YU!�2�bCY�S��a�F7�.�����썍���a��_��y�mp]~c*�jrm[��	e2�m@u݀`8Xg�%L��\�~N_������!w)�����|՜ysַ�������T,��6�=��o]׷��S._$������s�^gF ��j�D`�0�A6; �����g ��8�DBO�㖛���[?����֮]���'߯��ٲ�N�9/�/++�*//�D©���YR�t�$�Ӥ�&�"�����<���;w}�4��L&%{3�G�{�'�u͝7�s���?<���"�5. B?���׮U�;0a��ޟ��9�5���V4����DB�\X��xS�u���T:��+޲�C�`
�W��eƬ���ga����ǪU�J��G;�/gY7ڦ9�q����CX��nZ�d��=_x$�z?ۆ�oI���f.��NAcMm�iӦ��?�Ѝ7��?����qz���Z�zu�UOU~u�ڙ��'��o��BQ!b��A	A
�������� �������}�!
��A����o�u׽[��������ӕ��
�����Q��!vq���g���Ѓ}'1����m-�J��4�:Y�}1N������_~�nlK{q]%��P��El�ް������۰�2�/���z9g�**��6(*1Q���*H���nipl��)�sHX���0��ެ$2�*�4Λ�X���ƪ���?�Q��64�ڽ�}��5��5%��x:���X��E'7_�L��h����E/f��xO��kǙ/�ʙf��u�SM�SU]�\���[�N�;�vy[�b�Y�zu�СC5��b���������3+��*2NSI֎GsD$��!�B �@E4Ϛ	��FHZ$	}�W�92�3(�nx�{�㳟}��y��)q�]�ܾk����ӹf|�r�����\A��B}���ʞ�I-_�����)��\ē�&�N��&��Ͱt��O��{���3���S3B&�42YP3&�����X�|Q D��1	��!��(��*��X�<������?LZx����|顱j��r�ʊ��=׸�}��3V�f��I�t6��8+�����\F��| �D\OQD�5��ܱm+�]䳫����[�yZUծ���UUO/^����ɓ3W]uU�����]�~{����k:;/1��k5����ti�b��J+�DJL�̣�`�"`��!VWuS��\R���s�~���������w^��;���7����>��6l���������a���ϖey%�h�#�cE*>����u˭����[�ߕЈ�"��F������n��\���_}?���ړ���L�\4T�Vi�r]Q�����_�w]� mf!+p# )Y�~��5z;��6N[��WS�;�f����ɳ?����������nf�7�h�`�PE&�R�$��c�'h����ݐ���l�K���0�.���FdY����tcOEiž����ɓ'g���2�tj�޽ڦM�b��ۣ�vm��� -b�ϴ�l��Q��&�b�jD��ɠ�@�f�U">� HA&͘	��`��%q�Bax���Nmڿ�w׼�=��Ww�|˓G�����^�����#c�T[�&�nj��y8eeee���~�=�`KK��x��?� z�� �֮-����S�����<�\��Q�du,iB����A���.)��]Rd��t���vH��,����������M�����Ξ��06�c���o�/���v�������l�L&S��f��o��9~� �#��=�1'��ڱV�=+=�(��n�n.�K����]պ�{4U;�E��������7+**�\.�����<���GE�`g�v��@���c-��slۜ"s�u]h�9��K�c+�@w,�q���I*D��b��U):h!�h��RX��j`�0�L$aDbp2�������I�g���~��HnS�F`���_����e�oO&�!\cu	j�u熡�g���f�ҥK>��j�6��<!@�~��~��9��3��];�L��OI#�y��TeX��g-�P�1�*`;D�3�%]Jc6��+
�*�i9���@RT�1)�r�N'�P3s�o�.������Do��/��R�ƍ��_���v�F۶c���H�hA����l|�O�Ð����������?���{{g9�i�y¶�>U��4U�e�[h'�P�+
u��P(��4�6��B��i\�un��(�$��9�dL��,6l�T*%��$5���$F*3�L���z�uj,˪�k�U��u���8f��DG�v\0�Cص�VS�A@�4m�k:�&�{�P��P?m2L�=���X�8�Jtr��'-Z��i˖x��m7���׾v��^x�u�I^���FO��M�Er�`ˤ�>��O|g�y��?����b���[�L�������;ԑ�d%�)8��:jã�=�@¦/�LSD	�h�:f�g��9HN�!����S����|J��3�>��v�	�`l:�=���կ����dW�
�r��Vn. ����:u|ٖ+��Hؾ.�c�eo~"������0ގ����#�T�ٔe��T5�$)�V=�0Y&I�(�s�H ���w����m]S]۵��)�Ɉ���r�q� (IR�19�n 8�B�Ǡh2�2Y��H�s	�By@�j]����q��r h��J$jI	4L�����F#�ST�8��{�zj�O#��Fc�oqҟ����+���}��-�H�V��3
�ڱB�kk��ܴ�m�>}睟��'��v�H B/�ز%�m��	g�i�X�{���j8N\Ι��"��+X�!Ԁ
.x9&�y�11��*�8�7m;g��Kn�]S����efu�U�۳?�I��]���ٹw����U�l�r��DEQ� �&�v�D�/#��B�!��;�����`��W�CM|�S�o��;��q_3�1�.����9]�4�mP�q8��bW��l�<>���g��ֶk�"1I*Q|�v �p�P�Q(�� ����)�mj(K� XQ��r��x1X�
��,�e�}�`�?�._�m���Sķ&� ��#��z��g��4��Xo�g	�d0.�5��߻����W^�w�J��@�_ �9�Ț5e�7�4�s׾����Kt۝�ZfH�:�=����h�a�N���"�p���Zq��q�LS�[��|f�]j,��nZ��ͳg�on�cmmoY�	��9p`OEǾK���,f �QU��s�d2��p����sH�B��#[A��f��vQ`���k��9��W���~��'G2Gb�����kt�9nCE������Pۏb�9LD�{�[�,�?���[\F~���P*k��A��@$��rۆ�iC�Uz$���RPKJa��fz2�t����-���sÍ+vrж��-[�~���?~� P������AJJbh����|Ǘ���������_D�j��}�i�;:�"wfpQȲ"�l@5s^�;���-:��� (�G�^��*J�0���8�8gz֭�$�p�J8��\@~)�8aӄy3_�n��]��, Bi����c��ړ=��d��,涹�\����c�A$�|��Y��g}x�)*��V;�=���<�=� �<yc����/=,������$j ]pMW�'�\ �,��%O�G����Au0+��K�d���.WP�P*�: 1˅80�J
Dp>�=iH���Z�zI��H�2?ieׇZ�9g�U�dW��W���w�S���g��k�v��>I�,<Q���#�iz����G����/�X�����.� BC��k�����۸�Ս3�v��=52+��k%�2x:��BD�!,k�-[$ˈ���9s��PPX���@M:&K��	ǅ��T�i�k&O�P�ں�t����Ƥ�e�ʕ��G��w�n�8v�{N�6/7mk���F�u�m�c�~H$_�H�ǚ�[V3s�X�(2z!@���y�Fb��佘�{�< X㐖 s�K��r�G�pG�:6�Q�C@R@�|�)���@]�z*� �� q�AS�KӀA,�J�4\M���Z��B���F#p$1�!�W=��]��9�2�Lq�q4�b@ ��{�Ww�켗1V���H�s-��g<�����u5Uw��?� *��;�c B?�x��ِ�{}u[W���{���g��	�J]��a'���`7/E��Ow���&:0a���� 2,f�D�֌�@�k�̞�t�ZY�jݔ��7-�������-j�Yt��׃��l�Q�y���d&9��|��f3�2�΄�ꨎ�2�����	��M��eLT�E��=��'h#ڃ��0q0���.����7s9p���@7<8�l��rAd���o�����%	B9B.�M������kԼ�UMT� ��5��p��vfJ"?����)_<v���F����տ��Ͼ�jժ?g�"W�1�u.Z�=%��N�>둏~��;/��;!B?X��3aF|�޽u{�n��{���pⲐ�6���\���f~��d�5/�]�8���r���$`6nc8�K�UUԵ�ۖ5`�Ne��QU�oB۴g���W7�n�͞���Ä�m��b{�*���.�J[*����d׭���
�W% �	-l�Ơ�^���2>�9�e��Ex$�`u���ʢ��Y��Ǹ�_n�u�
� w9��\(�qՀ��AM0 (�� �.vE���}��>s`��I2�(p&	�AY��OL�n��U�D:�cu�����̙3�~���=�}��V\�&R#( 3TVV����0��G���=��+t]"�qr�pΕ�O<Q�kÆ�'������O�t*G�Qt7�K��E����-ȡ E@��5�*�Ta�TIYV!�ɂ�Ȑ�\A�&c���q��ש%���������ꛛ�زec�H�O�ʕ�ƺ�E�;;��'����iV�jrm��f�ζ�J`,θd8��,�Q۔�I;S��-��~�Z�h�#a�8<�2�%¥�p�P���6�6� �&)P��D�E�A�s(�E���d�2DMX�AM���* ��,bU��Cg(	?�tÊ���}��6��8�lٸq��/_��===���rj�)G"�'���T�x�g��O�^��S��Ѕ���5{w�n�9t��3���lvb ������� �eT�.4�E�Ʀ�Ԙ"z�{��(Ta (2�T�3E�s�+�.�[wӎ�kr8)G»�5�/UO����u������Ȗ&�utlw�=���şH*��Ie2��T��[�9��m;Å�,�m;v]tQ��q�qm�q8cgH��e��9��g̰b�%AI���1�%��I��YX�!�B��TU,%�M�}p��� 5�(�d�A.d`�<�����_r�W�?���(x�i�K�y��'���S$)�uݜ=w�3sf�� $����%9i������3���t=��Wܺ����}W�>��`Μs�r��R6aI�qE��O4zЊWf;���NoB��ؘ\�	9X���a�Wrf1f�,�/��.0�Y$�����p���P�ƞҺ֑�������_���	��i�I���)CCCJ.�S�ɤ��:!�J��L���r��8*�M��f�3A@�(z8����D�Ŏ!�����֫�-�C�Y�����j�B �����0����t�]	X(v$
�%�ߩ(}�i�o6}�C�.�^�����:|�p�K/���d"y->��&M:5s֌�����=c���M��� B�X]�[b��-��l�v�����R�i˩�-7����b������@@�ٳ����ђG�RT���1�"�rD|�K*d1�g[0b[ɜ,�ښ�O���k��VOj�^[?�;�\�,I$Rl�rԆ=/��+W��4���  IDATpX�t9Ø8��l��<x�xd�+�>plo��,��E������ΘH4�*�I��a��p!�2lV��i�m: +P#Q�j*��ў����%K�Ϥ�x��y��qq������[w��� ���I�&�8m�����a!���/���cx��=8�꫕�v��{��{�3�C9s��˕rǕD�c�.�q�`
&�Td�)��,Z�J�=�u,�o�'���w��mL���t�r-�@vlUΦ�3��r=&H��ЏE*j;��e�uu��"e�DEiE:RI����sYv�U'���r_"2p�he��=SO<������v��{�����:�갫��X��BX�K���H8�y�p�J]� �Y�q�2������[�X�5ﾱ�ih�E���3]u/�}��d*�n,�,--M�M�����Gc(I/B S��u)"гzu����m�x}���U��V�u+���.J�t��v�� ��#���E.Jҩc��ً"9�yt�c�]$�9�P����ʵ�+kV��i��.�&w�"�Ɇ����K�~,ZQ: ���PII:�g�lU�kl[U��H��\55�5[��f}���ض��ׇ��j�LR(��?I�W���M�M�sUZ6[�l7�I,RT%�Y����p��A+U����t�P�Z�0�!�̀!#&�� S5!�k:�#��ǶDZ[h�r�Iq^���[��=;v,ߴe�m�n*//����}s�θ5)o�������T�i���t��\ޱcϤ��'�����f9�+:\�0,� ��^�vGb�|p���jESEM;�9W��5�:��Gmy'_gb��6G�U �a�9Z��5�k�.V��-��#C`Ȓ �8N�v]�K����ȮĘ+�.;�s�]����ے����U�mWp� pM��궅����3�{/�������!ik�a�%m�e�)���Lpd.j����l{�� �J|DW(u�Ϸ\����]v�55y���E����P��/�����>������?�>c�݌�1+-`H�i�"@�^�s!�5�aCi��]eGw�^�����H�]��M�4�rK�4LC�<�~�[^�}s��$�Y�
v~c��Y@�A�f+�	d��r0$FT�Ru]$�����x$��cIV��E{��ߑN9��]a�KL�\�sL�C�8���%���t��������V��tU;�� �cQWH�"�K"��Z��N!3xM�8���+Ȇ�LZ��8�# �rE��I�NZ�dC��+�/�|�9�v���+~<<<4���Z[[;'�N�`mm����U�D�c��8:_�Vٗ�+?s�D�����鞁�͡�)ӮW-;���� �eÚ*\�H��F"T�R�D���z��)&���-��"�ZQ����v�O�U��k��s��;�������#1���қ��b<���A�ƌ�����\(��_X����#pl��X�D�5��Zs�������\-GU!)��t@������W<_�x~Y����� ���j�����oo�GI�*jjjxsS�&M���H���.���)�Ћyv�`l��A}��=5'�8s��u=G�_��\�;��[vم�o���Đ4���L�f���m,Y�5�mT�B��ȼ1}-cg"�F�f����w�G|��o�\�}?�羮繞��9�6�eT�4���������h��h}�{V���+Ȫ7D{湤4i�X�%�G���t�v�m_)�K�kĝ�rw����v���/�Q��W�Ǫ�;xspK�J}�j]�o�=�F|��Dw8��
ä�UH����	.�s�X]Tta�����ƽe�E��X�$0vDύo^�u<˹s{��(τp�I���ba�&�C��=pzq��#Ah��3��E�GFG���rÁ����/?�tӼm���^e��B�i�~7PN�i	&�s*��S��[���}������躺__$��m�O����D����1���B| G'�����Լ��j�ԈU�T-�5����d�o��`��ɯn��)P~ɦ��y�����y�A�;LQ.��F.(�إ�.&!���gݑ�m#��}�j���l �'O��q�HgJ�Y��4�)?���al����.&��.v�N_���>!4�^���I��'�
/B�[l���IjTc3[����MK���f�����d'�Q�
�)�Cܚ��?�=��	�N����E8��'�Vm�Oϐ�qO��xE��"+���dVC8��kB��o��D�i:g��̰��6j9�6�J��ٗ����^F��8��6mh�M�}���;�;�ۦy�X�2���F�w��ߋm����1�� �pa��q���CD��܆��F���)q��=�����go�����Za���ts}v����ɧ~���!�gEte��<MO9��k�0 ��1��,�q|�f�����������n)1�֘��Q�1Q�[Γ���Q�x�*��S�-�#�&)��WF�0]^�"S1�����=���v�Xu�Dݠ)�kn~������7VN�G"��B}G�/�Dq�]��X��9c`��m&�����غ��

�Ӷ�t���x����_
�z�><��	ɯ���3��oT��M��%���4ޏs�|>G54�^���ք(u�x~<-��s�{�jҙ����fa���Rbʒ�K��P/O��_,=kC����G��d��͜]]�i;�+`��j�-M�(T�P'�d�k-4�RR3m�\֥������چ���*)SBɒ��YنA�>V�}��|]�8���v"ּ4q���_+`�w�;X��Ղd
v6����G�Pf#�;\�	Đ�I$�]r�E[|yH�\��F���PQRY\y�[ߗVHcR�� =8��(+ݹ�{0Jp�OF?�4荁�N%wLsK��<n��}a+�H���|�	�/Oϰ5xR\�՟@���F��כ�'''_�Ɔ��r�=\{���1>���
U,Mm��̛�a5���0'�i){|<��a����V�-�,��Q��2���@�!r�9�
Dʑ�j��)��Fy�8a(�(OW�S��&
y�c��a9��Uo�i}�I�3��n�����^rz���:�$,�����w�a�V������3[�^�+�������y7�`F�V����lx��+v>���]��V�5��>&���\H�=���1�u���~�e%H@�b��L� R��ō�n�@�����x\U�����7�2:�(���dֲ���{�:B��sC,Ȍӗ��ɹ��JK	�V*�����>����3��g^`�f��5�mi�]qݦo/����Rii�u��D�����^�5�����+���/��.���2��QT����~�g}��U9�Vg�����i�z���qHI�*ldƃ�l8�ݳ�j�{��ݽ�R0j��[���7�7�Z<�Nؒ�55�qqT����.eV���s ����H/n�NBHb'ݎ;^uزWS��	��{(�I	�i��%%��9Y�����P���2�]���Wzv�/G~jU��֚G�R�X���@��,��Y����@�ڼ���U�飤�[�iĲY��$�ğ<e5dX�H�U���}p��=g�(D,��ߊ������gl;�j��{,F������� �0�& ���~�g��1�u ���py�q\f ʯ���?,L���e���L���b ���k�X ��4�J�:���8 ��w(X��s���0�E��;(�}�i%���~��?����	��>4/SP��0���q1��O�/{~��˞�S{VX)�}���� `X .���w�PK   :�-X�L�,� o� /   images/a0820d33-a834-4c8e-839c-8eeec59e25c5.pngl�s�%0�-zڶ�i۶��i{ڧm����m��}ڶ��}�֭���I�Vv*�T���ΎTV�F�Ǉ  H�2�  $  &�$�w��?�����f��  �J��{\t[�ٮ��<	�/�2�C��"G������C�@�Jb�*�ȱM'Mӽ�_&1�)�;dc��.0S�l�Q%ÆDE%�b�$g��?��=���W�����|潕x�)}���|})�;�ݺܺ���U�c�^����W��Xg��P�_h��1��8��q���/���F������Ai��������?VXdZ�����������u6���7���"��d��p�@�l-� ������9�r%,oM�?.L�)3�ͤh�L����!�H��iۜB�%|��D1�LH&I��e͑�qe��:�%�H{�%�W�Wz��ꙺ���**C�ɫ�~�T=wI-k��/7���Ì���e)?#)<_n+v�\n�j;�x������&����Z��~��mઑ)d��U��۝�И�ѳ�<-�x���]�hS]�-��J��zx>������T�H���K?�v��k=�{Up��p����S�����M�Ae�I5�ID���5
���4u�,h�G�uR)�?HQ˔O��<�n���4H.��l�����IbfZ �(4�R�*C]
��&2��*u��
x"3��M�o��}릊"_Xl����a�2����A������/]�/��M*Q����?���(I�WCD��� ���Ec�o��kr>�i�U��4��~Y��yެ�U�FCRE�S婱kI�_z:��k�mA]C=�\!�8o��mU��[�B�r9�Y�BQ:���	ċCT0�YJ�8�]�%f��f'��T+�j.B��A��h�q��-�ApL��Q�%c��d۬��@�7X�̈��D��e]\tp5���VխwV��+TdO���m��T�����0�N�=�4���4؄���bS�}R�ca����^��_[�:�V�_�:,�l������^��e��s��ڊ�#\Z�����{�Z�{��<�[����Ϯ�>�H��1�޸�Pf�d���S�R�-�ȱ�իhT'��� ���e�B�C���L�"��Ѧ
���2	��� �$	�XU��@guIץ$E�✒��*r�?��ֻ^�v�n�ȱ@B<�1�J=�� ���gn��)�Hq+��[RE"����q;A���w����O�YeT��n�5i�#�d�����{]���!>�� �v-�i�JP���F�BRH^��NTRDJ!��R[��<﮺�5�&����d1l��x"eq�2�iYK\}Rj���5*Eno��"����>�k$����2U�X�)�PY����m����#�OB��^���jUU��3������=�L��($�*+�����,�R���6a�7�9�b��/ӮG��"B�����ū\�v�z�-�Ӝ�q�4n�$���kMQ-�9��sz���V3�-%�ZjYE��1�A�kc�æ�:��Ovy��dko��N�#bP����1�>���+��	��?|�x���N���NeP�����u���4��c ��ף6�F����ݴ��+z =�%x���Y���L�а�+���^�\���G�0vЯE�1��`c����HP���2|�}NC����~g����� ���b��4�K������׵Z���[n��R���L��ETӗ��ЙN%���"8���u��t(�o�����7���J�}�����׊���p�8�]	M$�D�t҈&6ڰή`�#ިL#.����%�4���:�q����}�'E��d��qʜ��69�K�\�!�, :�6>O�?�|@��JGZCw�C�Ġvte��A5�C���v�����ۃ�W������������?#qW�{�]���>�[[�<բX���x7�ퟀ������t��؏�x�w�\�o��{O�S޾��w�(uϧ>Bv���6��`c�;8E)�N��Qɱ�X��}���OX377���,�Kn��zDZ-��P{&�aQ=�&6Zc/�c��q���9�Y��f�����_
��h�"������ۮ9�Pz���?L������V{WG�\�Kȗc�Ê�gc�aIdlS,H2��~�nw���v�a
$]�IJ���*yg�0F�j��p���=��lu5 ��������JA6;�-���$�ʵ�p,�,�b��&=���Z.�K�Z��*Ö�1��X+�Km�vRl砯`��Q5Îf�`�qY�5)�io9r�Mତ�>_�Z���N�D}�aC[�$���UÐ�M�͡��F�8G��[&sV��)lr� mJe�&-l��9I��b�ֺNV��]!�i�S�sml���%͚UY�չc/�L�b�lAos�9q�^s-E��MS9-�
X���i�0�U�	@<���6�d���L�s��F�{sŶ�i�tT�5��<>�"��V˲�Ȉ*M������Ql�^6&���0p�G,;m.��>EA����:�F��
����T'��������n��i�_�}nl�Ñ<�\�?�f��<��/54R�~�^ϴ<�P٘�Ud+���ũ�Y���q�۬Uw:^/�
�W���[^_�	_�=E����޽��|��L{�Ѝ�@U�R�J�BgQ�,1����f!�&��D�Y�h�F�MNc������;��������|F�&.#p�� �(*@X���0�a}��/y<i*�7�{>�z<�2gϜ9����&[�
./�B~��v[��T���`O�aac��H����R���$oHY~�(���#�뱈��i{�70`qrK�!��$��./bR�E��|����ndp$ؿˀi�����P�O{6@0+��(��iW�����x���D�w� 6�� �)��U�dl��e�c������_�F_��Ӆ|�gB�R�wx�@7�����Aϡ3����C��ځ"x��nE/�TҦ=%>Lf�X>��r�磍%9��F2F_�Cp��U4�zp�j~&�P	
peI-�^����ԑ�
B�����v����4�*��!��'�^*P�y{� @�8xxΤ?��ܷgMY8���v�G��?�����nyw���E2E/��p6ؖ��k�����D2�L��-��l�T\��6��3͙��g=��`Z�5cw��
[�<��pb��GB��?M�KaM�ڵ�@oeں�6s��\��EE^��V�:@�1��\T��òg'��v1�gt�d�m#eDx�>`h��k�;*l&����7�jL�LD#b��k��������ga�s�봘l�3��%z�U�`S��WSJu�_�&�F��F�q���{�'1��9k�/�����/K��}�y��?4E~��~J��ߵ\e.�E%:����r�W���։?���ڹ�2���v��N�-���g���?�V�gQ�.~QB��;9��ݎ���oUZ��
��8�� �<�g���!b�;����Qfq}�;�_n��w-�[	�9�r�&"�009ӂ�����~�	w
͐ma  @�vI�� ���+���1x��퍘M�������l��#"5��6�0����wj�H���ؾ��,Z?��}cF �P��qZ��Њ�]7����2����#�4-�?�!�WF"E|�S�f/���u�>$o���ieaZж� -[�ʸ�����D��l�@���F& �����Q��p��}P>�[���$�x�C.X��2;��96�N�
QQ�a��>�cpg��X:�a���W�d�XN�К]/#��/��:�>D��v�?y9�ZɋMsX��I"F�o��x@�e��\k'1uK�2��}		<������Y�x����:2� �p�JeG���s�<(=��a�!���a��΀�ߞ1��rGh#p������A��Ë\���\�d'&�b�OX���拳�ǓZG����J#�«r���©)W��X�?�<kQ��a+�V�U�m.u�"[a���p����UF,��/�;H��h�0��d��k�kAe�T+\˯�p�[�����,��<B�u<�՗Z�'�>������o���Մ��A��E��-�KG/�WA���$�K��~X��x)X����ʦơ`ϑϝ}x�Yc{��КZ Y�h�n�sE�҇s<�
�KU �
�D5����]#e�}�9#>5՜z<Wy��k5s�����ޯ]��u�Թ`�$��G%K�\QpO��!u�ִ��g��SA^�M�W��s�]���/[����~�wGs��^�=(�w(�+����R�)qP,�h���Z�͟�"�����
�٤�F�`��l�:�"8���lF��0	FP��7+�Y��>�[$̉��C���pJ���.`gF�R����n���s���l�|��]�u$��wt�6�ɘ+�NW�{ �|��߯�(?B��o��4L�<��;���͝��`�	 ��B��o`�-�V
�X�M!�oR,���$��D뤣,�5�_T�0����d���sy}�l�u.�>�'�Yd=��X��'��w�qШ�G�E?��L��
�}��4�Y�?�ά\�h	K��-���z�v�>pA+b�*H���n.�
l�F'�X�&.\�*��Yoo~�V���F�=?<�w3ǁ"0H��~�XR^t:��;��҅�$yc���Fn#�Q\,�~36c��k�n���\�H	� �ѡ3�1O:��W���ī�2�t䓒���V���K�b�� �ݮ [�t��������=N���4ʦ��'p�pw��&�+�}S� o���k����ɕ���܂��"e��!녻�і����P	�c�y�̐������,�:7��:{�O�ֽ�Ɯ5������L�~8JY�^�[��G��{ w\��7�ֵ�%�	 �_�w7�%.�y�ͽ�c�����W��f��n��V1(�o�|2$ʅ��M1�<���V�Q�v�.���>Ә�m;31��s<c��X�n���N{wE� �<3��TJw؎o*I��r�7sQ8
�]ߞ��B�/7���Nk�|�&����E�zߟ��r�.��E��Īb���a,_%g�Mh�ġ��JE��n�iϯ�Ks'�|Bx4$�������ml����J��$�ρk�l����ZT6�������k�Kg[�DBI��<=m�3SI���7�g��H����~h2��u�!7\��Ԃ�0qjY��X�̽��ɔ����EO�)�� �m�m�"��'�����,�;��)�Bބ���F =I��
}�,/?^TGh1*����"(Y~���˽�O���}�Z�xo��2A���=aO�=5����5l�m�}ƎZe-#kmS�3���'�ꀝ��d�� �5��,&��^j��5�@:5���f[�'
#	׶��0����T�!O�YUwe��y>��j�흩G ��4s�vY�F>p����������S�9���е#�An�bL h�9"�GR�`o�%%&ꇕ( �$i*Z�M�.H;H��B��7B��`��ӣ�U<%�"�WS0�A�d>k����X�Fs��D����z$!��LJG��@IL�9X*lU=xJa&0t�� 5+�tT�~_s�^�$�>��NUZ�q����Ӱ8��=�&�P������l�Y�/�H�Iy�:�i�� D���߁ف�Q�EVx&&*� �X�^�-�$sH'$i8˜99{�7�ɨ�����R�*�\C�(l��H*.�+�����e��1�	A�h/�S$΂,{��ޘ��|w@�э�̍���.D+�f�i,���+e��Α�X��ܸ��0嘶���to��v�v�`��AN"bVx�4}`��Or.���C��' �lú�5���QOGb)j2�
yN�ܨ����8�jB��j���̡�K�����s����C��e�^����1��L+���ؗ�澕a�w���gao�>L�kΩ�6^1:�
��cVRMA�5Q���x���5-z��𨿨,�j��՜x�)�G1I@��2>_�n=~ߖ��苷���/#�?�(#�&�r��|6��w]�4�w�܃~��О�.�KܮK�~�/g��hd�v	�*4��I���+T/Ȣg}�u��+U؜���a�=t�$�۲��MX�N��]M� ��A�H&F�0B��u�5K���6꽲96����xF��h&��>E�&�����f��N��c�l��t��a��r��������T�>RRҌvaHȣ�,��=�Ta�@���{2�#n���z�;�p�Q����'�Je6�XV��yC4���`�����~�|��3?�@i��k����I��WR;��`f>���f>��_Q_f�����_R���LNI�������ɕp��{���<�w����Ow���I��s��S���<�]��9�X�sh[�r�H8�6�[:�	G�U+C�mB/X����7j�puu,&�M��ʐ��x3%]���Ћ�^�f�r�� oS�T�D�|,(ٰ1�!r86Ҭ�1	'�4�N�g��r���҈Zj�!�^,,���[""�Pˇ� `�u,��61�����[и�5�����~Y*���Ime�'�B�߶\D��c�S��4xڜab��>b8G��l��j��&������e�#���6�tT�� y�aI(r�4�ۍ�g65�)dbS�;�>8qe�^������m�����~ 8^"^���>+�H7��/)0�Uy�˨��#\���:�D�щ�i�'F�C�ǿO� ��I6�!S9�O��T	zh�Ҝ+�m',;�q�,cCw��I�CC����@��7�L�tn�-��1����i���N;����D����]9��g� s{|3j��s����7��`瀱|C@���} ᮳�KW\\ܪ)�3`�nK2l�8M�\|b>�	%�R�&b�^��*����=���M��Ot�ʼ�n�(��Ƞc�.:�c2"v�L��#�Q;�!��`{a6FU���&;�tĪ�=�\�R����Q�﹕�7j�W��}C����� r�
L�F�(��v������z�7�.{�d["�%���I���6��y���m1�f�T��+�š�n�G��t���Nk��A��ټ� �r��MP���o�V����86X�Y��K�J����.�\
63��� �z�v��f<�Ƅ��ۏ$�|ΖK��US�F;����g(�#�^mz�J_i�E*����y��j�=�ژ&k^0#���X�u\��Lc��#�Z��o7�7wf����:�-8��B�B~X%~"��A��yΊ�/�"��8��{�ۋ��xO W�!	�ԑ�rϤ�s�SFu6R���b`x)W���ilT���V�c�c������A��޾��}�ߟBx'S
�Y�����Ǌy�ӿCx��*g�g���e���瞤��O���1&4p�m�r�}υ=ϯ�;��[W�O,U�K=>�_����l��V\�
�C.xG��5�H���s��㫻�n��%�0�H���ϋ�QD>�'���OB���`���}�b�޺�K��6U��<�I耒c��G\�o�\O�5��a�F��. w�#mL�����ݭ���(R�����V:Ȁ�.��ՠ���:c�d��8��ujȿQP8��t�6)�2+��S!,t}��c�Y��l��8�O�</84��X��m�z�z��W�?�9ݤPX�>�!/G"�$���}�ģ���^�y�1 B�B���Hn�NI5@5���aT�"p�)=�ǿ�G�������WK�f�l
S����|��y�T�����.�8+ C���M��c��#䰉��V�e��M�{���[�D�bC� ��+
KZg���H�S���%�3�b� ��XƐ{���߆��i��[�;��eÏ�@�=����/1��ՏQ2�N��Z����]���U2�;�D{M;=��	*KY-\.;�Gx��l��X������D�P�R���� ĨB��I��eø��y��f�j��p�	TNf�8:�O.�TP!ъ%�����z�2'��:������ľ�G���9�����B-�����>�a�Β�Q�N{o�_�mY�c9+�ư�PA��	$Q�-�tɀx =�Cb������Z�����g�����CǊ���L�9�#�O���^�O��|Ɍ�t�j{���m����8�]^���g���&z�u��!��HSƯ���G'��pv-�bqi�4�2�硫#PCP��)��ʘ#�Pf=k�����z�?	2Z��O�Z�d:�a��6ȱBf�NΓ'��P���)����@�5�O�p����|Ya�O�?�C*�xuLp��]{2^���UvN�}�[��A�pF�2r�E��y�4�0Ȭ�^<�%�BB��&��2=�і�앖Ҧ��%:��Y�aS\oo��Z�c���g��!\X[  ���3,:�{eK=�^�d�}j���Y��^�f!��?cL���*m}�B��O��l�`.v����O�1�
�"�H���j6������6���ԺԮ%2�-h�dI�A���%VM���`��a�����t4�VҎ��{ߐ3��oK�C��w�/�OC��n�?�&�w<N� ���lv|�E�v��^�BĻ��/��5x�DCl�!���$A��g+9�Ԡ�g�S���Wb��L���Y�v�5�7���<t���8w�¬
C�4��tG�GM
 ���bzP�JR_�Y���]�ˤ?$�o�2����%O�l���q��L{#]4���������ޕ�GI�����|�XpMg�z�^��k�u��r-k�/�'�q,�57��1�f���'�K"�V]0�ߙ=�n�KYRfG��Į���x͌��5M�K �e�C�K�g�Z���k�F1���+�{�׫?2a�W�\8ͨ�Y!�b��TcF)JadS��Cc��a��'��7r<n`�#=J��$؏�أ��K	��/8�b6 ~�?�|��n�ĵt����tY��������A��/��{���m�<j�5�I�tEpZ [��)T�o�����-1#]:U����_����Dm�C���7��t��i.?󼤙�)Q���+�~w�t�z�I?����U�.i��\:�o���v1?��d�[�m�� �5G�@�g�������ɭ+^�I��H�w?���;�y�$t	�ONR��X���j���=��)*��}�1���������5��C�����y�Q�!"�I�� VaL��C��OT���7�=&��~��yf�,�E˾>p��^�zyE�`�O�?C��'c"��P�q��A���,LCǇIq���ҳ��ic��#ݔt��t�_��93y�d�<g�[/�e��K8�ݳR��;V{��{v�Z���k���^(B�r���7���?S�_j�_��%d�#��q����#�<��|Sa�	�P�?��[B�5�a�E��~�ĽE鈚�6�;�I��b�̽��-��7?n�7!��<��`vI��۵E��]:FM1e��x&�>ϟ����������J�ϐ���2�aخ~~ɒv�P'���`zA^18�q���J�B�;Y0���1���6�Ȱ��{9-�%�k$;�sr*#��5�>KF��L�5?�|h�����	��ǃ��[�H��V��a%��h�-2Ō��߂����������C�+���i�8N0���e܀k|}C�Db�d<3�g�p<�Q+ I�� `�0bۧ}����A<�@��{t�8ࡔm>o��[@�5�9���_��^���}�=�Ad,\��	��l��d�����I�{���	�b����0|���e�|��.�}��*#7df�[*F���^�,7vӵ�������LV映A�,j~7IT��tX�$(B~TZ����Ƌ��9uǞ*ke���If�>��@�ҴUu��G&�PYR�Qw��]<j����	�����m���LC���7x�fk�u����8\������B�ݮ��kV��9L%�C6�<�=�;[��(_0�6��'|�E�"[q������C���ޯGLqM�*��B�/ �������gR��AJ��v!]�ɼ�	a��kn�Y@��SZ�JϑZ���� * "�Ӊ`00�j��'M��� '�~� ���?�6����6���6��t�sv�9'��	;+1��no�=��(�CUE�Gt	Irc�{~�ޝ$?�[X�zd�p��M�7e���u@�Ol�|�S�� ����U�����{8������gv�"y-���e�idT���h����`�M��{��[��F��W}9�,��@H��t����j׃��L!�Ǹ�F�%���pQ�L�/�n}H��<w�q-G�����[�4�7V>/:���z^�"`�k��z2�;�#�&Cn���q�%�����I��6�	�Y��;�c�!Z;������[$	�(��B�}��i��?Hm�x d�{�e����F�x��:膦D��;� z&I����Ƀk����~0�k�R��(�PV}���������i���d�@�������M(�M����4��_9���!4�Ş�t�#���dpȿ�����Z}�7�;:������FB,⟡
�~3�N�,a~gm*ZQ��_�����G/�$ѥ��:�v��F� X�0���a	-���H�T��<Pl}�F��b�1�M�h���z����|�Yek�M�Y�rm[�xNЃ~��uɲ��[I�� 6ۘ��1��T��kb���x����wtX2Z�y�}��bh���P�z�A���N���ӹnfrg��� ��g�Eʙo�Z�P3Tk:œ��[Rz2W��g5X���H�f,�'��f�(�d;*��5W��MG�{������箣+����ǇJl��͠?���wJ����u���?�7G������7>�Hq�Iv܉�Į�]� n=eb]�K������}Ut�w����<����|���;[���D��k/��V@�^����{:>���������y��
$����E������ �l�#�8C,
���t�p�����K�rQpS��<��! �Xi"��|n�<Ę�;d����s)���A�����)h6,Y�����$-
�%.<�*�4��)ę�t�$�Pw�ڌm�ｂQ��/Ɖ����tUbf��w��]�&�fܮ̦F��v���Wx^_�ǯ����^]�"��EcUA��#Q�8!ajj�-}���kޝ+�T��f禼��8���۟�.�����)�{ ��Ȟ�!��r��˰��������,�Ǔ�73)T?�:��E޸�):8��A]�SLy_�)��_;��y('E��wg�:�Jb�N=�A�*@�Ρsԕ�w��*	�d���Eύn�h�n��L�̏���^GC!�.���w�JY���\��h��K���Z#2�'�py��E���5���}1��g���cJ\d�?�0�1Z=`�g$V��|�~Pq�}x`��^�%���֢��=��S�P�v;O_���u��S�ʫY�Kw�
/��������w|����d4��W(�شV���5�ʭ�/ߔ��AǷr~���O*� �P�v~��7�Kz���D!t��H��z�z��8v~�tĕ=�¾;;�r%"�����ɟ�(�F�[�O����ԲB8]q��T���c�=3�!�Pb~�b�_�څuؓ<8(�d��&��o{ѿ�]�D`u��]��c�$U�9	B������?/W���P�U��OB9=NV@}���)�
=�|����]�<�q5��%�Ƕa�J,o�a��$��h�,���|�[�|o|��)��2�]�Z'���E��g��b��$�J��{�}�:�[�BWq!�55�H6����D��:P���3��)��6
� x���H�`B��<]0��/�կ����[Xfۭ.��;��ҝ�$��k}�r�n;�����~jXA�;��v�1V�"U���j������*��V�� ���A�8�9�	h%|@ã�O �5��Ob�4yMa鎦�=�3,EF�t3����w��e��iҨ�	k�!  �)�㡬,�+� ��r��� j��T(|lvN��=��E��l��5s���1��)�awE4���Fw��2YϫZ1gt���M���\/�
�9&��z%�W�gV�P�F���Y�>X�߀����
�����AZ�?i��z'�����en��Hf&�
�\f�M���i�U�$��*�/���|TF,�"$T�V�"�ڱOX�j"7_y�{,t(���z�J����?g����\�Au{!s	������+) #=Y�X%��=�佦�O��ջ�>#�GLGk:n_�:��z,�%񦲩7f=9$��HAOL���&��m4��-?�%�Gd�5x�oy�� X#�Z�>�n�y�C�h��*�<����8�0s��Ui2�j��z�c��R�?��a�z#���g�[g�l�+ �mLl�`h^lQ)�V,�x��eWp/F%����WxAD7��Y��ud�N�{�-����D�a�.�+;�ُ���u젃��>�ټ.󗉙�wo�E3����Î�9Kr~��q>�ݍ	x[7~��j}g}��BY���]��OW�։G��W�W+$����J58�4fK��N����ب�ɛ�J������Y�j��	����9g�u�Z�$�j���J��TT
2��5�3�-�ʤY�\�Z�n��n*�MF�Vx��Ul�qQ͌��uבc�K����qy�K�Vl7u~q���%I��E�%}��W>�hn�u4 7�j6I4�F����C���]���O�o��޳�:h^�oyK�oɎ�z���E_��$�/+�'���b�]�}�x���; L���.�]U^<��ǆO�{`Nb7��oc~O����;K<
�I�f<*M��u�;Ke7F�r���G:l�M[�$^��'�$>���`ɁTj�U�Yit?�lռ���|0�
�>8�-e
�	�xbA�� �S���W#i�;�"�� �,��� ����n�jH(0��^��y�=n��`Z�9n�`r8>�����[�c�W��L�nO�Gd�pH06`<4-Ȕ���8�/{*��ǀ%c}K9ܯ����j%���Ji�:�/X��G�4m���ABR)�_�U7Rþǜ}f�k)vz��p���3}�x�7�Zq�ew�U�c82�7�fy��$�;�M-.g�������jT5�ޖ\���|�,�2[��V�����dՎ�B�h(�ֻ$#�F����5���Љ�Ԕ��e��5_'�e�4�r�sĀt@�Mӏ��Rz+�Ty���^l�j=)��V�P3�%C�&؄��������d;��Z����yɼ|�6Yyz~i�����R}�U*�[}�xs1���C��e����`"�>v\��%}|%�2�@�6y��#A�Gѭ�2��2���4j���:�I�'�'�����J:�� �a�A�r�4m~�՞8��������9N|h�� ��1��Y�����g7a�sC�߿����c�Ѻ�X'|��R`#��{绖38����c���}��b��9�z�����,�2�!�?����R� �*�201�0�d� V��@��>oje�(��s�\�"��Px`�J�4C
\<koR����i$	����']a� � ��č���"|0���7v9��Xɮ�j���A���ɜX#͖�{4Jvz�5��y}��XM��fT�q�L!��z(�b�.k�����=.��V7�Țey�wr(N��ƒ/~�#3#{H�x��F�Z��ޖ�S�K�$T��Ş��t#n:��A@/$r���)�F�9�v���������2�,�j�f{Id������Km"K�r�:m�Wѓ�"_�!���W��ӊ�����=0\��@��*�r脗"�����4;I�L�P��\|��fь�6N���7j��%�ɨĕ6��N7�Z��rYWE㘹d�dTwgښݸ$.W�'L����o�A��2��0�_L���E�֠c��Z�B�B�W�@��y��F	4��>���|{�ҝ*����X2�P�����,oY��PSI&M'��_�Y�Ww
�r�VGhk�U5��B�ߖ���)4�ja�݅S(olKc V@1J�<���ZRS?��+	s����Gޚ`���u�Z�Npbx`�Zs�ȨezcEc�c�0�|�����kJ�q>�X�=b~b�Y4�:Q੊>�q��~a\k��Qc���u?'ga�|�c��5i��qLj�����V��U��`nJ�Ҳ)r��X�@\���f�L-�l���+,0�Nr��|o���������|�ǎcY�*i�	f{(�
g�KQ��O@�IsxQ��nYw&���]�mჅp�d"�Sl�C�W�Ǻ�0�8Q�-��g�^�GZ7�!�M�UXi}��`Vq�6�!(?;�eʣXyc�	t�/�X!�r0�u���g>����o�� }ɓ��ްSG���:����	� h�eH�k�c�6��2lkRɡb(k�5�,�ᬾ��,l�Ϝ������D��^�&��l՝x�y��>9D��J|ӘT���r �Ƃ��̽�[�}:Ӝ��7���F�� D�A-[[��K
ʈ ���}q����%�9c�ׅ��2� ~p?ʺ6�G�) ���o�V0Ӭz��P;�q�/���O'�C}p�09��8)��R�܎��n�]0�=��|įF�}-�C�"����4���.�Q~�{Z�D�m�i��>2�v���CS����i�g%�*��(<�M�&��@}�@�B)H9��l
�9���S�l��\1��F�Q0*	y9Xlr�χ������Qbx�y w��Ve�l��
'&�E�������Y�fYF"aR�?:��� �4	\��'>]���y���!����oTՒ�':���y�|���ݡ�"]�C��T����U>� �]��Y��^O�2`W���s�k~��Ӫ��w�7��0�v'*&L�m�<,�tb�<�O*�h�$�i�X�{�#'�d��/��ig�<j��Z_1x��Ǻ�����
<t�Y�RK	�
�B����F4%���z3��a��	o�y�r��6d�O®1s$Oy�R$�_���7*�����$�<�%O5<���+�ϛ���J�_�V'��5��#ϴ�qcޫ��d}�2�X��XT�f=R,���A��0��6����<iƱ_�+�T��(����{��"��	��䤂�ʨt���2��#�{pz�����A2Z��Z��`�G�
*��2�2���%�s�a@d����p���Li�!��A�71��U8ր������
�����i�p(��?k�e��D�@wSRRѸ擫e�qH^H�Y�m���o�c��[��y�����Zw*^]���ت �Q�ЪJ�3�SX�q~*����O���E���[oz�X�����h��'�$Ȑ��e�[f��PSr�����2����"S��Cf���]���ە����b]�PO�!Sm���ڑS}��L�=D��qAs��5��5��ɔ�9��3����,=n�ٟh�����k�@`l�gR���wh���?�Ǖ������l�>��ާ�<Ⴏ�.T�����I!���3:s$욆�iA���TD��ʾ�{�Ӆj�9������"q�M��ͽ�B�۔p�,��8�sw*MO~��a!9ES����p�t:P6��� >@Lm�pAY�=&�Zft���# �k�(J�E`n��x%g�K����Bbd�Y�FjLԘBj���T�U���0�Ǎ�$vSX#ƃ�ݔ���ҜȘF����M�;�z3?�>��G����'����Ҍ���b����`��?f		��ܟS[�;d��U��^��4�VՖ�D��$57#�-;vy�x�k���;����+٘��O��훧��h�8>9xp-r eLvm&�f��=����0�!���狞K���TO�<�WY��mQ�6-�9��Y6����X�^�������U%'�9�{!� ��%�`z��Rf�r�
�|��� &���n���\ �]�D�%��Z� ,P���(�*!q�
��(�r�x��:�'�^��܉Z�4!:����[#DD��e�6�}��O�
�Yf�����f�lUl��:j�f��jTrt�Ҩa��$�Y����,u�JF���_T���<����7�n^�3���B��@����3B��.�;r�V�B��c�Z��'R�%�'瓬�]����!n���g�	R o������lP�E��e�rF�
m �f�)��X���YX�%Փ���%txp@�1IF.�0��0�LQ�=(p�,���p����O��C횔�~��a��A�c��u�R0���-�f:^�X������LJ� c�>^�+Z�b�s*z	�EB�;��֭�N��dlx:�� ��ƖlB�m�y�����:�s<����3/c��w�d���2���oX/d\��>�/�c��~�DQ�Qǘ�����=9[�v�b��Y�8�y�:״!�B�8R"s���1���xko�� ܷ�졨w���d-|�_W��r��}qA�C�<���}���v<�P3�W)C����y��k�^��$ԅI ]�4���6�i�Ϲ^�ĺp2$6Iz�0��1�6�8�26P��H��/ �(����(����3Ħ���HӔD�n��AA�~ϝ��Rw]8O���^:��Iyө�u��\�Ѱ�Ӣ���!����콡���Θ-��NbM弡�����3OPC-�kz��-���O��{wsoq�(w�b�E�k�m�D6�3�!V��#O�t�8�lc��DD�Бr1䉶�q�A�P�Tڵe��^���_~�;?�����x����z�	��/?��������#�{0�8M�,�lب��Nǡh���Y ӂ�E���ل�\������7���ȉ��1��gEHӂ�J�z9=���B�����Α�V���sJ�$�¤]���X���9/TX�1��
y���D1R�ETk�>�т��4	�b�uz=q̙{!�(^�<F���V�����j�7|G��u��껰�{7;W����~A�@޼��4xm�nehB�+8�U��C���V�`i���o��yس���&]�����i
+��N��
qv$9>�	��b�Y��cZ�!K�bJmY�1g#���bB�w_����來S۔)�Â�\�J׮^��W}��I��r���o�bt�� �.�B[w_bm�k���\<I$r`} �] ) ky�2�$"=��\t2u�Kr{�b B l ��k�DD��Kp�z~̇M X�%U�#�D��|��-	��p� ��X�B���)�q(r��Sl�A�!�;�\�J���.�-^��YTP��˃�`H�8椀^!@]Ѝ~�U��26d4i�^@����˸�.��8�	y��EپZ��K?wǺ�ܓ�@@
�3җr�F gh;�R�dV�Gq�]��!�u|�0/Ej��0}t����Լ�(�����;�~��䞥_@6���b���i���1tC%�\���C��X��_d)�����Ue� m�P9������%Q�X�qbX�|"<b��4q0>�W&��g�k�΁[ק�%�c�GQ�Po4�b8b�N3m ��Y>�/J6�s!����Dn�g�K��"&����9�׶r��A/�(�t��C���V-o��`8B�w쏘�0�ixwB��-���g��d��}��`�	�q<� �Ή��ᾏ�Ր9�|�X��~jѰ�B�V!.{�����1�I!���Z��1���5d� θa���9�ܣ�Ϥ��q�3������'��H� O K�T��h��d�>;?|:t����F!��׆��nz��_A�~۷�w������|�*��4%S5��0��IK ��G�s��|!P�8�.��CT�9U�	�2�i�/]<CgϞ�5������SO��{4��TS� ���:��ݑ��BZ���1Xk@�00?�} ��4�Q���3����0�3�ktv{����q�4�s�%���9Z�q�]����e�;��8f N{{{t��u~��ic}�F�u��$���R�"�ƨ���tN_x�+�ȓ���/?M7v�6���Q���؛C����@��)��k=�Dا���(�x�-���5���4ۿ���������}�G?����~_rB�7>�����>�u�`��E
F0�^�R��Ȋ��ؒ��O������ɕs:�%�=��M���t� �v&d���iʋ>Q��M�1q��S7���������JS�Q9� =xR�bb�6����`��8,~��Vm��[���A*�f��"\�U���7���l��+&	h}HQ�'���F�u-7��hi�2�D�TX�|��T��e`2��Ӱ^�D�8���A{���	4ZRQd4��c2!���nx���ɲ�� ��~)T#�?�g�1����{���Ƶ��{�:YΌ�?OZV<�T�'��T���c�������s��g���[�Ԍ6�<K��=�A�/���h@�h@O|�Iz���|�H�� ��(�CZ�Y����.H���s+���%p��	������ґ2Po`�v\z�dd���
��bߝZ�����p��B0F0����)��Z�ER����mC�b���Ĝ�;YZ�;��EB�$!H�xK�{�1���S�lyo��B��N�]�]�=[�N�/��v�r�� 0�CPê��|�-�	B�J��ȧ$v�-Xw��t=1|� �ʀ�:��~�G ���v%Z/FTOy�#]����1��O�d˒k�����$�br0k���Gbb�Cpr>�G�Kλ�O�ɨۉ��cl��͒g��}��ҶB��״]�B���>�O6i��3K���l.@�d#������.��C �)����n\y��	���7b_M^\��ڐ���i�1�!a�&��Lx��f%��:�Lh:��Y �_K��~�T��Y�A��s�=�Ȁ�/!>
/6t�������Dx!k��Yxލ�i^!yDNk#::�gC
s �}��W�&&/ �a>�D�	P�*�����4���� x2H�����<��&�n��D���q\��e�s6�=�뺱	=�!�8X�CF)I�,k�����?q�R'�P�8�2W�X�� ���_^}�?)�"���1��oK8Ѵ�OPB�a��4eq��c���5M���aoH�.�[<K�{�k��s[��D������?�ǟ}�667�-���iNv�lr�x$J�jN\U��fo@�V������}��O����҅�b�[D���g���)z��}ڙ֔�=�)���U�9$�>�/H��!�����/h��Ҵ>�Vv~Dq[��SCz�+�w��Az�+�;�l�3-�ᆐ5�	����iw��n�i�`�IM@�ٻWW���G�nޠ[;{,??s�:w�Z���E`�7iP�TD��c���.>?DѻG5=��ez��k��S���2�KJ��T!&�G�K��c=��� Y�L�F�x�<`�PY��
��vB������t��������G�r�/���o��#o��_��?{�~c���x��cR���^�
�kG�-��re�$���)�㜴�i)���<H�ַ�9�:@��9sn��P�%)M�g�x�>�[��ݱ&�SKY���"���q6!L��:~q!�B6^, ���@�?�H���6XU!MLR& \iªy���`b�\�8����k6��E}��;�ã]^�Ξ9��݃��eEA�ۧi^���@7n��x��8M��O֣�����o� h[�= zl^�ꭒX-���$d�g�����V Vd�(K&X ��zt��5�y�:�ءvQzw����D� ��S�z����d�,^���nHT;e�,T�56���i��s�������Ӿ0�&f�G�����V���=	z��C>��%�fbs�ݿ0���v,����y%�P��),�b�|1O�.�Y��e��V��u��,2>��Y����S�.���ĐG^��m��,�!K�Xq���Q����K� �ˠU�J���/�z�s	���c�ޅ ������Ɏ#cT���?��dł�c�)@��y��%0Q4�́��6�����w�{=��6��^9�[C��6��9	��9��\�s�c��J�Y��*k��޵�{}����%'I��gm���S�a	���['����`�$AH��� (������B
� k㾉F��X�y�ܐa#p��	�������x疯BI��5���y�vk�E�N�>́�oث��f� /쇸o�s������ߣ[7whr�1B
 G�u�m�Bb$��4�Gi���2��I���s�"�tb��钨{O������hkk��#RR�p> �G@���km퓍��a��]JJ찞�y��p�s&0��{8��ձ��K�����G��x-���W��X /X�!s%ǅD��hg����
`w�A/�``2�rގ���������Pl��^���>v���1.�ťd(�+@�@ X����h"A
H�v�Ջ�C�1u��!}�;���tn�8F��=�,��?�i����[��V�ѿ�#t�sH��$FQ`N����*J��"����=��c�g�gt��e�#K���|�w��wn1��b�DtX��<J?��E�<u�����Krr:�iYq%n��:����U̗�!c4o��܌6��x����7Лx%���Ktv�g�:<Z���!���'�'��_y��\�Ee�Т	� nHR�v�⢵T�Yc�b��%cSQ�*z�;�F���ҝw^����
?��3C=�8�٣�ӓWn2�r0��yCM�Qel0#���J�OP�+��'ƇWq ��=s�NomSY���gh�}�-�����_~�������4�_��%���o�]?��?�3G�{஻��͂k x�T5U���,x�,,�����v�%�QJ�`�־~���oz#}������4�xNY"�d!@ʶÊ�w?�}�c���)^��Fl�iLI���eI~��/>l�q�"*�Mܖ�� ��w�1��Ŕ����vT���CS�T�3j�9-JE��"EiQ?˩���&��.?�4]��<M�3f}���>E�.\���5"h^[:8���tΕ-5�MQF�l̓	�6*X��b�e�Zq{�,� *p):��=! `Ɇ_����3���s��7Xp�{��v�
5�Sjf�wq�}��,C�&��DtA�2S
�A@?�^�1/�� ዘ�Մ�.�2G��@���w���u��sj`������ <yò-�ʎ�̋.=�M㹄B~F--��! 'A�H�����! P>� �9��� Bֽ��,-�'�ju=B>�L�%w��r���t�������aC��R�O ���!�N�J.�G�1?��/&�A��٩��ϗ��;�u���sK�mG;��ba��_~W��� U0$6H�'D͒؅�� �,#8Q)Y��������4�l�.��N�� +�c1
 �s���Jb�}���{�uw�.=)ᠥGF,���LAÒM,�a(P&������ϫ�[� y���C��g*>V<8ȟ/�k�XQe.t���&	��(	R B ـx� =A�w�.��I��E���!��l��� �m�`dr�τ���h6�����⥔���-Nz���A�.��� �&��0R�:t�'��ɓ�"-��Bk���[3��_̽wp��}.���q:@ {�$J�dI�-7Wٱ�8�'Nb�nO6�7s���&���l�Ȗ��b�rdY��e�.Rb'A��~pz/;��/ �z����� �9����W��3%�+Hnn1�z!��,�J"�Չx"���>}	G�a(��fQ0�@XA�5�S�jq��҃ό��>vdjJx(}M���ܜ
~�]pݲ��`��F-o m/�i\�f��:h^�nx*�1�e�C�7x���z][�0ӠQc�]7�����R�v�'a��z-��1�T�A$4���'i�	Ѳ��6ձ8�t���q*ڎ�ug�Cys����l�L~v\-�ߺ��ʢ
���!7��g����+b��9>!B�Uq��;8��>�;T��66�4����
u�{���w���C�����F�J,(�G�4c6��w�5k�?�h9;1�'o�u ݝ	����qގ-HE�z��
5 �����,��އq���hh����F�A��D0J/�P�V�?A���j�r�zmO�������g�F�ٲ�{��c��X���xo<���yL�;���9u/���&~��A��JھA��c���z�e��j��J��R.�Pȃի��ߕ����صmvn۬d>�c.SÑ�)�|�8^:|���#]n>Ԫ��H���\�!��F�T��5v{L�)~f��b�]�������cx��>wr�ͫ���?�����%����~��S4ٽ��.Þ� �m �EǶa�(�Ј�Ag����_��o��v�`ƺ	\�w/nz������d�j7Z���#�-��|?~�����t"ڱ�vPYr$F�e���J&�Z���wgpl;�X0�7�%��zٴ�k��3P!�nToPP>OS�lJd�*�Ky�i�3�j�vD#X5؋��AU�'Ξ���3�Uʘ��B���AG�
�NmP�)���/���>��"�3 (�IY�6Qap��iA����A�LE��ʩ�O~�����:��h���F-g	BDU�zM	I?t[�C?{gN���TC5_D�R7	�HS&�pd�`��0��-2yLTf� ����"`��B�9�q�6z֯¾��BW��STj�fL@Ņj$}:���*V~��n�K�6lۊv��/K\���`忣C��5�3q��A�99���M$\����@�܆��w���,	z�Lje��3��=��ҿ2�w$Y��J¯�^��mp��� ֋wE}�D�ARܳ]	���__y�+�s�VT�Wv����wH3!�J�\���%K�Yj��G<�圸���Dp)p'I>��w���W�	C�\�Kq����
������ݼ[�3�_9�~���Dj�/�7V����0kz�ߛ��T��5���XQ�zg�b��������GBPk�K�X	u	�f�J~�6-[��9,8�;����;Z��9���=}M�L�T`���VӘ�Y��@�T�db�+HB��xϪ>��[���"��-r0e��: U|�5�̷�֫"!N�&�4h�(�N�ҕD�B�
��_�������P�����^%�8;�B"١����G3�VP��Z��:�w!o��`H<�� <j|�2��)ty��*igF�?mV��!X�Ph������N��V�%La��\��"n��!|g��g&��?��v�0�`��E(�)�2��+;�,�1	 $��J���AC�V[�A�V�Pzz�B�\D�8ʵ�&��2���)@����NO>����ќ�9�W�B�xN�O&����I�;����O���r����0��������}���җ�� �}�O�{����3�����/�1�u��o�f�-4˸-YV��J�ɩAމ�3���-�5WQ(Vqzb���\�����`:SF��17Wk�C8�D��}d��j �i"�i�VȠU+#�c��Q�{ׅ�x�6��I!�"m���Gq��)=6������ؙ�N�2�2�'�?�z�\PJ'��f�Ĺ�j![.�ή �lIpnӜ�PO�Y�>�Ԛ�d�'�YF�[�Po{/؍�����۷�w���86Y����ŷ���I�gȗ�1a���6�6E9_�A�
�|��R�H�\}�mۂ�x��_��3;���Oܶ��_��2#��?��+����O�x�������7�r޽w-�?d�A���d2W����?�o��C4�1��Q����w]��/��R!��%��5IZr0���`�<��!��'ϡ��@$>���ļ �=d!C<�\f�$�	.c�Ȉ��nA�"�����6(�3��MUD�A�� qg�2���E��yx<54*%�s������n�F��<~���̴���BI�~2���Bv�"%�B��w�w���I
����"    IDATIt!O"�ę��#��cl��2mJ��r	�ad[FUK�9�47T���Ȫ	�h�E,�i1���c'�xf�lA�87n)1�'i��]�r:\,֒�/�
��L��觀�I�j��!��2-%׽�twczvJ$��AW�R�$.�ҹ<��Ym���Z֮����j�w*��j����0��k����X\1Xq��*��	�J�y8oo�sfxo�p)�/��گ�נ/�T!^��k_�<\U���b��̱D�^�����_x:�A#��5@l��.�|��_�A}DE��Ļ�w�7ᷫD��!Pm��/uf�ׂd��,���s���(��2�{}�,��x�qj��\��;��g�y���H�.����I��^�ڴ�_�ߓ������R���������		��U�Z�ad�n�~�Z���+;z�?���r�l6��N�����B~��G\ �J(?�zK]��"3�g���t�����O���'I��Ƌ|-�ZS��]<gR����X@����ٌ��B:��ܜȓ]�$�����Eg��+�1r�X���L�AX�G{�l�+�f��B�N��<f�&�P�B� ��5�C����4f�^\D1�C J�ZL :�{�9�@�ܢ�� 1!0P[�rF�K{�t����b�H�֭�b�KϿ�N�:V|��5�&�$[����!�k(`:�ũZ/� �	r�� K
Z���T�*�%����4��"�,�ݝ��	����H��HX�=����l�F_�b�S���F0G�&P����gǁI ����u	�zo�������P�;r 4��Š!�2��3�\�ʏ�k��d���S�]<���.+ׁ�"jo�<A��,�GN���(#�(᢭[���W12���8�u�w1�0��/���̧�k�J�*�&� �bx� �(fq��YD"1���Q����5�F	�)fpz�,�?���������<*M/�7nC��>�"'�e8�V0�J�:�h�Y) �:B�*J�9�$�سs>���{�ZtG��r�N�A%���O<�7^ۏ|��b��Z˃�� �y70$�/	��xP�V�-Qn�Q�7��V4��z�ZEB�H}!�,B��'�@:�Wǫ�(#�[�h�0�ߍm�7�]W^����80����๗_�Ͼ�����}���C�/��/���<2��y�y�z��� ���ء��?:�{��W���+���}����������o���Sg���n� .8ob�&bl�0��ߐv���|z��\�?�����q4�>����q��c�7O��f���*\(�p�(�*�c�ď|	�FB�h�C@��!�Y�7�gS�1���nx�2A��m���Oh����׊���Z�~o>V��y��i,��^��%�C�F��A?�*[����<�3�L��02|�ή�� �x��Qk�-�7�@(��?G,օ��at�E+�o(���H�n�W�h����B�<7nHt����d'�洕Jă�H�'�M�Q����dB��ݭgƄ`�3/��-��h�=eR�C���['�@ΰ&!X
nY!vf1V���R]b��hPثUT��o�����u���Y�,�����S.y&�j��ʠr)�uxj�q\�O���`�ݟ}}zg���
fx	�j1+���[ɺ�%�qm��|�ex-N��(3(����b-�g�m����%׽�\E��c*Ӂ%<�6S�I���۪�Z�"׵�kc+�.! ���Ҭ'��Z�T��Q���D�ni���V��4�lR��r�<+�U��ߙ���ǲ����0�<^��!���<
7s~�iu�)1`�O�� �V�F�w�k�N��D�����G0�����Z� H&�	��XԘ=;_̼p�� ^��s��C^+���m����I-Ã��ip�vM(R5sS��k�$�J*���I�f��	���K�� �s�^.�����"����(�"	�;ܼ��#���診�l�O��xƣ�'�.qf����W����Mɟ���b:���Uv�\�������:�q�z�^�U���p����oFc*�*/�7L2q(,�b7	vy���(gq��+IpI<��n�����|r��8���/ޑT��{&ć"����3|�/�f]�+U�R�ཻ3��7!=;�g�yF/
hpn��G9#�@4F�ZV"���$�����$��Pz�)8��U}��W�[�v�S�|&��ǜI]*���8t!��Q����(�s��!��GЙLi��;�	�013��^��N�����l!I��&����AK֧���
|��;;�u����A(���c�/�P*V$R���£<X(���IX]�^��1���	*d]���7�=�5�>2 �W�?3���t�pZ*El�W��q���8|�4��ޝ8t�0.��|�S�Ɩ��xk�1<��#"�_w�5�������O�M��}Wc�y;13��$��؝��S��Co������019�3��X̔���h��(��hE:�
DPg"f�°��"�&��ڕ�ߺ��&\�qF��-,�6?�o��Zf�G�P̗04�����'(�҅�d��:8,2�d�T����͢P-#W� S(`!��\6��LN�B�!S�r��l��\�"�"qd�9u��s��
�����p��ׁ�G�$��N��o��_��|�'�SB�Z��&U�
3��ٿٍ�2W�#������,��g/ٶ�/>wӥ���K���g������ppͺukї�#�E*�@2G4��UCW"���A��c.��/���'O!��B��@.W�ڑ�8��]�Ivjc-䲠c#�]8��|��S�q�C���'܏���u~��V�)�F��M��i��Zx����C�Bh�.T������R1�z��Z��z)_%����|!���
�b!��&P+g�!�0�QՁ�W^y	��4��L�%�����#�CzqYV�8���K>�����5��$:�=0����m��0�v��
&�"��͕)�CK&����P�++v��X�!P27e��
*�p�e0�M���/��7_z���ޫV�9���*�
��X���A���LB�T2T�
6��ÊR�K��
�``�(n��&D�b�MσF��G]e�\m�^��v�ו�ʯ��ː�Q@f��qwPSq[V����8/%���d������3�)֌�k�I���,���P0�7s���@����Y4��8930�O���*��� 4�%r���6 Jx<�:�+�"]�hx���DQ
�X��#�x�ҽ]�9�R�"�3�?�C�P2h�[���e�;q��Hu���]'��u��͆���ф��b��`O?�-��u���Y�y`�`a;Kl'9(SR��͍�G�5߶�X��6�v~�޼��
�M������e����C���I�ҐMH<m���9��;s�I�3
i. �j[����μ�R�1�� VKɧMd9^"��(1Au���.e���(���"9I+(`�^K�w�1��7LZō"&���A�#�;�c�9t����i�`>^���T6/�J�V���5I���z�T��j4|~]��':0;5�.1�><b��*��F�C`�_�D�TCde|��4*U�6i6F_{��"޶|m�y�~3�$�l��S�a��N�ԅB�K7�~�u/	%cXI���'W����(�Z�*1�}MNN��-H$"�م��!�T��L��Պ ,�/={M
�@��ȢS�^����P�����Т
��-��?�52dANґ�:Z��: ����p��{�g�Vv'Ѫ���;2dW����D�v��k�rUr�)
z��(�S��������VG��]�v����E11�ų���?��8:D:Ht"_��� ��㔙��j ��VDe|��}�����@*��!�~�~dE��s���p_�g�M���	��P��1cµ��d��=��Bѐ)Z"�#�0����l��Hg��� y��?u�zE��/����}�Jg�ϟ�9�{��Ţ��oæ�k��/������?�
��[���[��?}���w�N�q�m���[oUru��I�b�Y3*��'p��	A����R�3�b��C�&��������x�	�Y���m��9�PEg���m��k�e�0PΠ�Y@{!���$r��"
/��W)^X��xB2�{�L�#��v�����B蘩Ri?*���U�(��(q�PF��Ʊ�q���~8~���D"]��y��_g��5Q(����[�����`����*f�|�����+G�&P��P��W*�MO%��LY�%4�Z�[m��]H_�q�/?��������zu��C�}���>67����v� �ѶT���Z"��VB?�����|�3�Huw!�J��<3�`ڱ-�Ѭs�-+ �?TB������@�cH�Cd�S�2\t�:<M���!?H�����9s��k6��Zt'�ڐ*�4rS(��\ *y�B^$��o+Ȩkf�,�!��d�H�O�^�jE�l�d�b	_�Rֽ�C��F���`�_����DiV%�w�D��#X�q.�{9�mہBӃ�s3Ȗ*hQS�c�*�_p!TM{2�ep�GA�,�me�k��t��N����_�th6�a��~:�&����o%~ߙx�j�H������θ@�U|M{�%"��`������RBp�-7!�����������^�eq-���AȚJ������vMlB������T�J��]7��V#-��7 �=?��*��Xղ�2��T��}3�bgȨo���#�J��l��Ir0<V&]�@d,�t�c����$0�#MG���*oL,t!\��|5�pQ'>�ڬ�lF��FU-{����� VA�#�Ѝ�Au��S �b޶��;� ����J8���~�� ���Z��2��`��u7�ҬgU�9^L���P6n�����~T �P�.�^b������U��2,A�ͭ�lӡ��Ս�<p�flAK���6����I�)s�H3������r��3�3a�oeB��v@��Ѩ���2�% �1(�d`��$��n%LB;�VV|���6	����O�@�! n�td�cI�-�Q�	[S8��h}i-؎�2*�_��sNΔ/W�dy���[35��`�<�X(
Z�f	�X}=��1Д�G�9U���K����:H��G6�E�X��S�呞�E>�E�#)�p�3��U�"�P��/r���VrA\"� ^xoJ/��.�c�g��q�@���8������Ln�߇���I����Z�H��78 &|f�F]I�f	j8^�ȱ���uV)��B>/֬��/^{�eL��1�k��NX$Ԗ�f�HTѮ��،���^\q�&�l�Ƨk�i�z���@`-����9eJ^.�g�yw���YY�O�;j٨��'i]�E�����?�2����8<>�H��`TYo�K�5{1;V���F��������7��2�i�;ͺf�`~nOC�7��B�Y���Jf���"Dl�3���pU���_Yj�^l�ǟ�#�>�#i~����-7}�>�
u;�&���a۶mX�n�{�E��?�?*��Ƨ�w��c�?�o�q��������jt����:!�`!Q�!�0�Ο�?�<<����'x�WQ���O����ƫ�9��QDeq�VW�ކO�|.޹�F	�����<�
:�~���Dc����1/��j�e��m(v�!&�"i�}$�ý����ڰ�ܖt/�+�ް�;�����4�x�U�]�����MT|��J	��s�>}�2�1\��qۭ7`Ϯu�xK����^9x�h
�ҥ
�ݨ�����1Z%߁�̞:jS�nW�����n�������#��ï]���~��3��j�Q�@��T�I�X؃����^�wm�&wZ*1��8��q;\����ԼA��L%�	A"C<F/`�<��|�G����E8�J	A��l��4ʁ����w����J��uL�{������+hיT4Ѭ�[�F97�v��-h�R���"��J��[D">�c�L��[jʕ�Yͬ�5[�S� 2���g9t$ސ�Y��ڑf�{�a9'3�+�Z@�6���v�ً-;� �H��2��%��X��$ܶ�2���!H	X]t�o�1�����E�"T��N�b&��'N��+�#I�:�1���؂�Ky.�2n��&n��Z��KL%��Q�&A����:�o��T33�tc�T���7���/+��L��`=���0��j:-�������d魐���Vvڴ�Q��!/�N�B���3ash�."���	�2�5��d�,J
��ŐNB�C&4Kɞ��aaF
�D�RW�kMs#���IV2�0dp���ҬWѕ�𴦅nA4��Ye�aƉ����)׺�L.���v�,I�-w�J��׳5�!)�����-CԖaΗ�[+�o��(�g ea7K�dU=˷K��@�ڎs�v�%O0r�L�Y�6	2��m
.).���t1�<��t����t�򚨁Oe*cH
�8�R��ΑU&����2o[�3�y[�+\�uEe��f��L:8�Y!6��Ց�\3/�DMV�U�5�-Wp��F��5���i�b�=��HH^<C̼�uj�9E*;&@����,��b7j��M�������kv�:�b F1V�	��z�:�
����#K��٬�WJt!.���bf✤�׎���uk�>�\3�$���P���|=�C���B�X?�ISٰ<\���\wN���>�s��U.�07=���iq����.�����l� �P��H���,�*9Ƅ�r��1�7 ���c������t�?+ۂ���Kч�|��Y=M\y�����n�e�C��:/Y�[�k��f9�5��|H����-�����ߪ� ��� ��)I�۵I��X��WO�������W�������_���;`j�bA����}�6���b$e�\����<�*�
�'�5ǋs_?o!�=����w��ּ
*&��kr=(	["se�z�g[pōOfp���kwܩ��?�">�������R/7��8�5�n�3�?���D�q|��Ob��]x����;��1��cþ}�FwWR0p���v� F�x9i�ZφJ��ߞǽ?|S�|�n��^T5��_�h�sH۸x�z|�kq��;�Աx���Shf3TH�H�B�X0)�U�Z�JE�$�sMG�q��uͽb�B0�h�'J�,����ɇJU�H�D1��1�^,�#�x��i�J#Wc���o-�XT,P.,b׎M��-7��W�E2
<���{��819�L�^xC�u����a��>xCDoTD�Jhff�m^����=�{߾}oo�-��o��W�!��^�����f���e�4X��P+���o����>tûq�17>��o�y;w`͚5p1��ӧ΢Zm"O��d��x4�v�Y-����Ӈ����l-o���	�=�1���:2����=L5�A8�xe��J�ê�D�'hPzn3�c�ΟC�݁v�vٙI�|�%��b>�ba�RA_K� ���KRTGO�D��>��bk�/����l���i�l������ڋ�T�p{�B�<ۭ,�%1zޅص�2$�EV�Y� �/"ޑ����r]lZ}iI���	�������Ot���r.�srܜ<{s��A��JMʖ͛�9`����	BV�
)P��9oڊ�	�����Z����5���Ϣ���#�����!�gq	��C��w\�rh���XrKfpo	�a��Ӽ�$�DUR�nW`�MU��4-{%Fݶ�e�D�Z�vl]�<�B�_6�!K5{]D�8H�Q0נ`_�|��8�����^����B6�AC�s�u��8N��t'\�k K���t/�ī�U2���5�K��)7�v�\;����DR��5(r`�6�C��V+�I7�YZ·�Vf��������籙P���R;P&0\�x��4�A����N+���C[9��)w�T��z�1 5�����    IDAT�ָH����d�u'����b-Ui��ej���r��f&���|�����Ӷ���sLE��n���bCX_n���
�����̾�=�R!�|�~$Ti37�N��`-Ͻ��d��p}��t�h�5�.�8s�-u(�I��l3XRUۨ��9� *@տ�:IX�{�p�x0xf �qd��u����;�1_���s:�]���,��:	�60!i��Q�Ǜ�`��&=�?��%�[�o�1���3�2�R&j�~	r	�k��%����(Q5WĩS���f"�?�
�7n@G*�t6c�&c���֒�bR���3G��Ǒ�19~Zɀq�6��*蒫�"
�^kH��Y/#�8��+���o~�\�szha���T���<���4m`���e��@�L]{�LQM��oQ����}��mE ���-�݁B�{��¿�y7�{m?��$"������_���:%t�|��O�W]��}��غ������"z��Ou��J�	[�w]_��.Z�n����&�v���"�l�UM��U'��������G����u%3_��qۭ�U��z^䌁q>���q�]w!�H�c���܁g�}߸�N�9|����믕QeB��Atv&���i!��h��ٶ���8�{��:>��'��T��� ȳ���6�*�q������4Z���<�����,�QX��3��nkr���NXL��$�ٮW�*dr�۔4��4�;����4�PYT��ĺ�ѳqH����px*�W������<�m��$��]�ɟ97���p�V���[pյ�� ��ٓ815�v8��B�&]�)y�H�>�4Z5ʙP^,^u��/^��?��o<���� �}_��v�z�;����^��,j���
�D#�c�;��p5�ٹ'�<���86oۊ�n��*��~���uشi�	b0���H9Ħ�՞k���(�}ߋH���'���	�&~BnĐ���a�sS�;�!&įS���*����*��8��3'09~��<Ъ!��!4�]�O�XXB��E�VDoO
Ѱ`;̠�\|	�٣��?D�R���H)Q��h�ݡ����ge�a�K������1P,�
��i��.ր`���u�E�y�%Ȕ*���7���#��\mV�e�`�kӴ���R�ȯq���`=�^�b��)���їH��ͣ\,b����8urLwڔY���V�]�@1M�̸�M�X Kҵ�����
z7�ƍ�����ŜƓ�(iH��WXr*�>�r0m�M�7��`86 Y�t�A��p���,��@[�J�pӖ@�Pђ7I�d ��]�z����[	�=(������%I�G�ƃT$TV���%2��Ms�4���{z-�[��\b���V_��;e�e��J��+�%F,��yZ<+��̸2�p���I;v�P�$9�䏁�8&�6c��t
�������8G���-Mpv�l�$�w,)�Sֵ�`�9,���]���=&rp�LŪr!50O����ɱ|f�1�6�$�h;�-� 3@f�j�TPl��1�|^&@1္fC UR�"��7�ҥ��k�r�f�ױ���W�o���8^�Y���j	��R��ƵՌ9����C�y]u���[#T�`*��א�]�ŭ�L�nI����j=߇��*2�`jX���;t���3�)-u
;�/��$OL�L�����_�� �f�2'�g��c���A���b��/T2���vE)Bx8'	%b0� �&�م4�S���� �Xyg�J_YI93�\��ĸnq�"�V*:��;���:7�J=]�K�M��҇�l�Jy��EB_�������V�8~�8Ξ�T�BO�u�ף��W�b����N�M�PdSA7E�#hˠ2½������z��ob�M"����TV��F�|�VQ���ĭ�₍�d�.̹NOL�E��h\�L3��[���-���{��[�d�f::���lAG��qGV��K$B����b/�qO>�"N��F�ƛ��9��hI-��x1�c�{p�%{�q݈����Y� ���in�N�=����O�+�`G��1A��ipn�+,?��6�G��� b�{I���b������q�=��|�w>�+.�Lq�$�QtĢ�N>���p��D�>��ؼy3�x�	�˿|]	���8.�p7�Eͧ��Y�)���,��G�`����	)��O_=4���y ��?��/*�-�_�b!OGz�}{��.�h��gQMg�.�� ��C�vҾu����x�D��Eaw�|�tFIǉj`��>H^6�F��̹ �'�0��<^��J�E�p �nt��El�Z4�]H�|x��$�}�M�9>�s�"��I�}4 � ��Q;�����#زm=h����/�Ǐ�S�22�M/j� |�*������,�B��J>Oq��o��/>�����J��_.����'_}���~��-�?D�,���|N-}�
1�����	�����;p��q<���l���!e�?���;y;w���/ޫ�/�b��i�2S���X{���y�jI�{���iA��K8N _����$_V��˙,�t�:�C��F9����4
����;����y��5�bn��,��W�f�jQ�W_��4:2�v�������_��~�"�Tj^��q)�Y�W��yF�ITT���2��&��T�%�H�j��� j���ـ=�^��[v`&[D��@�ڄ/G0�6��������tu�+�V�M��3�[��J��N 7�FG'g�073k\���F�w.bf.r%���pMA�	�yo�d���0�>���l�x���4�A��Krft��B1��q|9�#��%;���`	+� k)X֢3;�g^c��|�¦jf!Ive��v� ��iC���� ~����5�H��y����n8B�����l3�,KRTG��\%R�����E�b�q�S��A^l5O|�d�׼�U�w$	�΀q 5��. fE�����@M�V�M��i�s��Dݭws��u@:���zNrrt�4q�5���بJ��J��W9�I�����;��C&q2��|�$���V?��?&�Z@K��%�}
n9�L�m�u���,��5�ƕ4M�O�p���#h���@]�&�A�!a`L���J��3�GH�_Lt%�h 5����re��r�YL�8�uг�ʄ�ٲZ�+����2$oY�W�c�^�"�d��o�7抦+�D�A�a+~����{ɀ���Z�Cbp�E����%�9gڭ��E�-�Z��T-�D-�-�%�zf� �q](U:3=-��t]�j�~���dD����>�7�ȡ�UgF?_�������Y�_h�y0���J���N�F��2�Cuu�Q���8��-���g1=7����p����ST�r}DR����+��*�R�Pa��'O`�̸$7�z���~�}J���DF	�<|��2ػ{+>���ʋ�#�B��+��_<�?�3d���]�c���X���7�3�\	g�F�#��ML����H ���OglGGJ�q�K._�B.�*�<_��EL�g�h�JTd@�D�X@ Boo?������ٹ�� Z�<֮Į��4w��[�Ց#���q	���l�ZX�bw�	�(>+)�5e�f`�AT�U��:J�%��z�vh �׎`hU��ګ�~��e|��㟿�m�Z�_��?�����1����2�ڹs'.ۻ�H�<�4z�!͍�ƓO=���###x��އ��^=t�������� fffp��1���P��]���oņkPn ���~�<�Г8>6�)}%x��J��
�}�^����"l��'���P�PFu1�]�g�aanV��J��&�����1�5Р�x:�������URvމ�`�6�L9P��Lg%ǌJ\���=���"ܳ
��UH�ـv2��3s��z�%�Y@��T?�&��J�ʅ9\s�.�Ƨ?�-�m��l��)<��a,�}H���x�:DyS&%�*�^.�k�F�
j���˶}鲿��7~�:~��|�G�S��g`���0ғ��YG1�I��k��������ә����`&�X�v�R%��{�ǩSgq��Waυ{uP��EL"C$�/�d����w?�\-����J��k�
�~�i�����;n�����
XUxZU<ĕ�P��`~�ʙ��'P�͢]��4' x�����Uf#T^i��ҷu�F���|�׭!���ڵ����/���"�F(���E�D`f�VI��_���n�i��Y��F-[�m���n���VP%~� |1�ۄ��}-��^d*u����~DS=��Ƹ�V�]����\|��x"��#��cqa�r�BQ�!蚥�������@A���
T�[  �9�E���
{"���xQMm[��?x#b]���[�k�j�j\*=���4*�8|�r�pڢ*��p��@�q��� �*U�8c=(;Y3K:���
�S�Q j!TQ"t�e�>��Y��j#LHxi�����d�FL���n�%�1�v]S�3w`����dX��;��S++�Rlj����O��E�);n�ȧ��:�q�������������1
b����Ʈ�<���wMS�3I!CF�_*�;�=�Q���$Dz/M:3V��0)�	����ov�̼���4�5�(J�aBOB�W�53F��e%E�OZ�������޴���o8��7^�:>46��R�:�ۦ2�H���=b㍳����{�"����򐴿,�ʤ^�DI+�,�[�e*0�5�X�XFn���|�0�|ZO̳�z���	��r$(�5�9��q��5�:r��b����٩k����h��.$��5�ﳤr�]2��k���pȯj(�K���L��~�s���O��ՙ����s����Z*����@oo��)�T��p~��b'�IL��S��o�5[�\k��Brε�v&��ަ.���{a����@	Yp1����Թ����{��r�q�|Z��7J삁)���#f]��Q��R����^�u�p��~��ҋ�Dp�����׋��8z���h&���"Y,��/^+��g�|��U{�C����o|���}��,w��hĈô[��X}5�K�i,V��c����!MD#���-��U�)t';�����WG���9�:3.߆��U�P��3��Ű�k��YuRXt$8M`frS���7b�M��<���sҥOuu���Cx��7p�ܔ<�z��DE)�\.�䧠�ʞ%�1Q�QY��r�:Ĭs_��k/���u����ޏ�^wS����������@�� ���S�_�/>�<��>L��UW]���������S�q��Dc�޽�d=����o �m�&���3gp��a%�?3�s����'0;7�����~�38o�6�����ϼ�W����YJ,b,����n����lH�4�3��O�!��U��\X���4ʥ�ᇶ���C��DWG(�Q�d��kv6'�Z�P�`��L�ǂ�1��1�-�:�斗>G>��X(ew���x
�~t�[�Ъ~�#1<s�z�����ɳ����	`��)�3c���>n��m(6��^}�?��fJ�T�(����\
uL�bT�O���6Q�?��t�?��y_��#��z�C����W�!��x���z������÷} �F{Ů��I.6:����q.�cH]W>hW��]���Ӹz�u8＝�X�)W�c;�CWi{���p���a�G�sTrج��EI� ����UvV��n�̨k�<��,�R�Gf�,��T��(-N�V���>�*<͊�Y���S�TT���^TC�y�Vlڸ^U$��ذq�|�i��������yD;�$q�/�u��d
�`D�kW��&�D(׆\э۪�a�<6:���]�����=�a�y�ETI�(6�H��B$�R��V�T��L��M�ٔ.��p@����TK%ɷu�b8}�0N=!'�v�h�7�l��`��a̉o�Lpf0�GkTvX54�!I�5J��Ї`��M���� �bfaVs��j�p��.*!`��%��GWS��?�
w�&�w	-S��B�x����-��b��m�s�<)��0�j������-m4��LB@�G�8��JH��R�~��eV��aBm�n<�l���s�t���eN��u��i��y�LP˟�Y���J�I2���!����z��BlTlx�.蕴�%�

�6e��:�	tww
�0unF�:O���@��V��3.�:�g�劬�>�:�ҏg"nȶ�NyI�٪���
���{`����Ӓ��0жr�L��y�?��hҗ�2�$�R֒��ȅUەR feu?��sD�9�
u��<Q��J��$�T=�z<��YUeM��`�
9�>�O�pwXc��%>�D2�	��,ɫڠQ��%\!1s�&�������NV�KV�;v~���&6�Sj:�ـRN2T2g�����ʃRu�ҵ�j��U2�������g��0%�	G�(����3j>�4o�4k43�]E���ӫ�K��P�T���Ic^[��x��<�5țb`])��	g�:��o�ǚ�k�#f:���@��s�%��;�da�]pI�SR����XH�a	�)ؙ�f~��n�4~�Ҫ�6jǳ��Y̩*�jd{��QB@YI�v��w0)
��"��r��0��	���x���T���]�a��*�;�cG��D(@�L�,v)X�$j��.ڵ��qͥ;�!@�%�����q���Ȥ.�WƔժ:[�$�I>l&�{��	��6mڄ���j,�ϡVXDw'��Wc��(��T�e2p��qIx���o �Q��)��@0��e1��_*U�Q-�0v��z�5|�C��ګ/E49J�`IA��������#�}�lٶMEV֙̜�B&��|wɹKh�G)a��m�ڊ_���I�k���}�b�P��O�}��lNyhjf���G�ڷ�����տ�k����'��?�1榦q�7�K�Et���V���A��E�V�U�\!���i^?�wzf�<�({�	$S=��>�իG���?��O=��c��j����i���9�Zq������?�ʘ;vD݁��Bu����E�i�3�H=����)rS��E(ͧQL�ѪVA�'��*{�$Kp�o!E�������&8X��`>�mb�u�E\�y���GD,���ѷm+<}8��a���\o����c�(T<�T�8|�E�������+h�x�W�!8q.�l#�\��"�_�X�8Y���5R��j(�'�n���{w�Zu���������c���W\�/���݆-�0\�٘�ŦQ-\��&�4�v��q ��N��{��Թ9\z����Ke��:��d�����7�����^��2�`k�]�P���rW$��"X�6~WY��"ul�S�� ={
��g�eQ�L����t-�iVU.��$�7�U�;:���f�n��:lߺo��*f�&��1s]��s:�z������ÿ@"�'�P$�\�dZ�0�a|�R�7V��̢`U��!vho^j�տ�?
�t���b��~�^��k6+�],���E ���aݶ��8��L�T�W�oL�
1�ԋ�j` �N��ēx�����d�O$,��0���˶��եo1�u]�[m�#AaQ����2���Xr� ����s�E8�0�s��j�졂Zu��1Ն�P�E�����S`Zւì8,���$=�*C��$z	��l�J���΍9�I�ɑ�M���v	MP{���!X
7�b6�d �l����r�r�*��ꄢ`H�`�bQB5�ë����EB�t�h#�]��4��:􅩧�[k׍����T����,j�*t~��Ãr�4R�jUt�m��ݬ��M��744���6�^x�����b�3��Y� յ�Le*b�?��{��'��|m��%OG��B^�cQB��H�;�*�    IDAT��1=;g�R@cC�N�'J�2�T�'�S�8�kv�,��c�D(@*�!����I%�D�[�!Ke��䰼�WX�+ԡ e���Tu���J����z�s��Ԥ�\�Ŵs�6
�� ¡$;����y 9Knd1ZUS&Ԥ$�uW�S��]1&��Uu���be��Q�,�=��¢QNa��j����J�}����I�ϫₓ��ڪ H�*���Kn:�"�«j>[ε�	�YP$����H(�R� S*v��0IfL/춗]戂u�5�b��w��d��K�?	��p3(pZ&�TJA1�R��.�tE�R�Pt&~^��}t�z�gV5�� Y�➃�s� �noֺh�����DJp �]1�0�Tl�Ȭoǘ��g@�P�4a���23=���oٲE��=3΂��Ĭ�pɟ�/��2��ǋ���C���H<���:;P.�8��B��\B�t��$̋\v��$vnY�?���㚽��A�D(�K����<�ؓ&R�Yo(�̂�6ދ�^���ܸ.��Q�X�z5.�{6�[����O>���	�iui��T�!���̴L�z���7�X"����r�%�htdH{gz!�`~��Y]Knq=])��u�p�9��fҒ��yw��1�g2��ʫq�%#�	%q��aLNLH@��+X��lm6���kC�L��
�܆�DJ� ��峨W�ش���ć�ћ�^R8R�5;���s7�}��X�a����L���{?y��s%��}�����o�+�I.���Ԫn�?�X���,�p~�hB�7c v3yj��,���^����i���?|���Pg �G�E�҂��@w4 #��n�W]��F��)�seDZ~��U�J��<�p$V��#&(rL;�����jTG���1���&l0���0�>ST$얜'#A�������8�KDX�x����8�jU������n��=��MJ$~��?ro�D�Mi����������?������s�A��b��|��
P>v �j��n�KA��
�g��\�������z%��۾����~�gϿ��7���y����&��d(j���D ۷��/�G�VA:���'�씋���?�3����s�X��b-���<��I�u�k�ʒ�1O0j������Ȁ�%�9�P��#J<=I�^�e�s��Ο���	,Μ���G��`�B�2�P�k��R�A[�H2���E{�Ǧ��%pj���E�H7nٌ��!�ݰ}�Cx��G��܏l�s��$��:N�9+Vn�ܜy�<��o�FpblL�O��"�6P)T	���uË�?�Vۏ�t��l�u�nۅ�JS]�v �*!U:�,,A��VR���C��#/rh��GY�dq��0s����$	�b�B|�$�9��r:`�y��+���97.r(�/[ ����O~{�� s�N��R�"���_U�
��E�l3�0������@S�kw��!4VR���%iϺ���N�$� ���U���ʜ$��h�ٜLK
��6%���ؠ���[��b6����X؏D$����(+��(U*�6�|����
�*��]���i8���>��̼<0(=����ֵ��}=qaw����аEY�FGW���KL:�Az!�r��B��R�*;w����2tnL3Bk*<X�v5v��.�ӫ��,c$J���(�
:8Ox0* �T��11�c��ɷ��[����ЮT�C��E�,������ ���qr�,�9B���M卡>7p�j] Eȑr2>��U�a�Ĭ���ݝ"�ML��R/��vp`Ͷ3�i���њT�D��뙖[�&d$&��/[QG�I�Z�'H*Eժ�U��1�oV+�HF��I�Gϖ��<�=���IP07�N��E�²D���++��Qs���th2	c�Q7]
�m|-�!<�:%��h�ZHD��U����I��ڣ챗�"?��e�U��p��~�$�k
sU����Wa�谔�H��»��e�-���C�;/옄�q��[ց���*j)hq�ۺ�=�5�G�o0�`���e�E%h�I�<��r���-�,�e�űfw��Tg���20�&���s�b�����@�(��Q9QşpD������ʰ�$X�4u�Fy��/��܁���AP�	H��>��@�#KsP�Ѻ���`��.$+��Z���R�;r� �:(rf*n���1�.sS�ٰ�ş�P1���Ů�k�'_�,��h�|~�D����w����ѧ�E��X�}B�^y�Ed�V1�>gu�B!�Z�͛7j�P���s<��A=v�Sf^�BH$S*4P�	g�d���mD��� �&},:��fm�C�:11v���\��(	�M
f�#��g+q��=�^MD���p����ȐG뻯�G?����81�R��3�f>��	t$ztمY���X?܅�~�#����Wr�N����,��|�;ߓ��W��㑟�?���t���+���oG<��;�1��$�a��ܓ��T��vr���<yRs��/���*%���x������;zә�e*��b��5��V[�
�p���a�ӏ��1D�E��'ʗ�g���r>Oǂ��b��WJC��	�3y�g��)�@��f��_u#��-x|5|�Z���,'L�ZA���S,��	��CD(�¢T�@:cq4�~���ѱf5:7nBǎݘ-6p�/�GO���/�@���Nc�����?�S9�����Cc(y¨y��7�����m"��Ga�j���@����k�������_����s���O��}�կF:���@jEx���$��kcˆ~�x�ؾe=�="�ٚիq��kQ*��o}�'q�W��/��	��#��BްI}��y`?�Q��=��������omB��7{[�%���ڵ<fϝ���q���d�Ъ�ѮЬ���6s4�l.�̸xDuv%�aݨZ����Vadd[�n����A�a��c�LϤ��K/���lQ�c@S3�:�x0����X��}��>;�*1ߗ�Z�m:;:��w��=*�������v\���}-�� ��Uԩ8I��,�:t�5U.��M%"�bRA �K�wavG�Gaj�%7���2�2 1�e���.�u0��gd�\�����9��C��F� D<����} ��=���ɹ"��?;��tFcvd:gM��w�0�|�:7\����V�}��)S�3� �Ã=X7܅T�A��HPr�M��պ6��+�r������@;���>�ZmUg֮]�M�Q-���Gܚ�u&�HD"�c�rU�Īa�#��q���LLby�.�Nn��T���<�D�Ġ҃U�������Q/Z�r�B�*�Ц�x$��e��U��t&�!���T��z|^BŖ	ܵfMJ_�u���ۉ�k�d��@I�,�[�OgEl\Hg�>G�q3D��Y^@�NV�9/�&�֮����Hă(�2�V��û��mp��4&&�U�����,M~�F�GJ���5�ke���p }���09^\L��kadt5��V�ٳ�16v
�si��\��*/'�\��+Ф�q�@�&���nqK�v��Vfi�G��J#}��ӝ@�`J�,� �����#c�x��֚d8���̀�R+[�X���d��K"N�_*b\{I�/W�(��̽g�\�y.�t��s��f0`� QIQ�L�"eYT��lKZY��ڵ�U�]׭����]_�V����"� �"�$r � �L��=�s���}ޯ�]���u�0�����{��IV.� Zt�!�/����m�0�߇d<���%qo�� Gf$s%�5�!�9��sU	��`�h��/]D5ή�K�,�w ���B�	�t��
.���p8&��
ϝ�A�&Y$)�u74;�Zڳ�z*�'���$�B�T�U������J&���w��!�Ic��s���kU�4��p\��EATl��}54Ԓ~��(D$_�5dc7KC��Dr
��^eq��Vm� �����M���m��׎��ݡ��u�Fץq��4y���p�D����-��������N�b�͇\�ҁ�MdMKQd�B:����R������y���yRBd]43��QM�2j�h�L�K�v�n�W>�Gؿk*��2R������o��7Ԍ�-[�������\D�(b�~yyY
���hmk�s�� +�I��pv�m��hnk�u��ōX��)�0s��hW��9�K�*/H(����~ШȠ�3�s)�Z�5���P_�3o�@CH�[~N��������%9Ft���@t��d��J�-z�;\H��.�#M�l� �@:FO������ć6�J�e�[^Y���+��g?GߦA|��_q����ӟ��/_FOOFGF��"G��!24�����!9�`���uhQ��x==p�;�GF_o?X",�%���W��ˇ���A��NX�������ܷ��-H��a�d`�d蓋r&�X"xt�Pd��������byjH�Q�d��03�{�܋bW]��Ӆ�n��� w�MP�l�j�D���V��d$�Ǆ�h��kZ��5`�;�����k���k'1.��sG�������f*[4!�� E�Mkh����Κ����[$Փ���х�;w}�s���ߩ������_����g��������i�f�Sď&��:�ݵ���^�w�������~���w�S����$~��"MattFG�˂U�TпX�T�Yp��,~��5�'u�� *&]�#d�G�!k���G�fE�����*<N;����E�M^Cb}Fn���|0�bAZ.f%g�v.�pJ+�:8�*�MmF���𹐈Ep`�<����*_���d�+R�8t7^�4^}�(���$��O왬�N���L����_��y�P��"��b��H��C��v��y����}��ܴ��TN��Mf]&��w�6��ʄ`�E%�r��
�ܺC��K�K�y�<̹,L���?�k\��hK�Ŝ����NC ԏz�S��u�_Ra��E�BJ9����k��<��|�c�l�#����F,	��i���#*����)�\��k�U�:��ZCP�����R����*R`QOUk��}�h
:`5U�r�t�/K��F��*"_&��
�ׅtXX�brvs+a�x;�����,�`)�:]3����H ��TL���*�(05��+WǱN���E�Y��2E'��r��n̈́��.l���ce��l�ܼ�"}�Ȇ��L&u[�̩rNb�p&2E\�1�p�3�j�T,�$����@_o|n;�.+l��5�=!��R
�SX^Y���"l��b?g�;A`����"��.�N���ׁ��f�4Y�P���s��l�t��lX�Hcni�k��'��X_QDbJ��!�#�Ci��s����q:��s*�	���;<.y�t���X,#��E$3IA1ı��Z!������./JU6�7������h4f)��N�\W�\;F��u����I�i6]E\h]�L��e�������k��p����w;�U�ky�\$�O�l�"�em-�L�M}4i�����l.���¶���6�c�L�B�$����r8�l��\��dI� �[��x�:��D�A-��L��NWR��݆m�G�ب!�_���KcB��:�K��,���01yK(՚�0]gQ��eF9/�P����f^�e���&�Z������q�8� b�����(���r%�Kf�p��3R<���s765I�µ�Be������3��z�!�8��-*��:=�_�kNtwL�Q	�k��5� _��ªU)Z� ���3|�l��0]�5�-Sj���h�˿_�&�!P�*�&�L#��9_���/cq�PkC� ��]"�|=
E� [PT<3ѩB
�T��Ɨ?�	��5���gAR�����������݉w��طg�����B�H�����	�(��x�'&o�
�uyϤ}੧�mtb�8.^������`�犡V���2���
AJJ#C�<�C.��p��D��5f�r]�@@ht�2�	R�L29�,�ɍc8�m����yvzN��x��r,h�I��q��9]�N�Ϗ;����8�V���3�r�z��=��>���5�(����~����_�����~��-�F8y�8�]�&���V�K��$-��tʱ��:����+Q����4��y�&�V����x�G��ׅ\�6v/���{�5��1%[��5;:�n<z`���#�G>��Rf�DT�v��@��]��')ƚ:ݨ�눐��JC+QL%`���$���m�@�Wj��u��HA�*$u�%⏢���d-�۫��
��-ҊH%ͺZA�fC��V�7#���7����qu1��A�R���	f�j�t�h
��4vR-IC�K`�U�7��k�w����F������Ums��_<t��ߘ]~���G�����UD�7�xػs�{����p��	���!���~��H�3x��aww�`����j�Fm`�C�-N\Z�O_���u�4��-E�t�r�Ň²�n�n�X�M�_���e�(��82�%hU�?(��Ş���9���v�Ae�_
�m[�����n��s��1:,!,"c��2xE���k�y�K+R���!������0{kJ���lA
���u�9{KK��L�ŋ?�vz�'Dw�)�A^�F�*;�B�@��6<���زc���"(W���D*�d:]�6-p{=*�����j�`azs�7�d(�0�U�5FQ*!�Q��]��'+�ޱn��I�$:�bLꫢPʠ��N���_�,|MA�l�����A6Oh�<_�D�b3.شw��5_���5(�uשh�ת���dUZ�Z P�ǜ�_m�V��Vty���$����S���i=��=#F�$r%��n����:Ƨ�qk~U`F
"}^7��[�:�T�W�D~�M���$�,X0,:" �.anv/�!�(��IQC�I��*!y�j�.���ϋ��F465���#�M���%Q�C@�䄓���N�+:A���;�)���q�/E����; HW&�hGmM�����"6x��9���,���ǡ�Wo��ʵG�(U5�+�X�B����J�A,6]�h ॰��n�ϫ?����x�h��٥5,�EK��>d�öM�(f�*!��2%��o�uu �w��q
���Te(W���5@����łJ��5L�ܢQʊ;����G8�ĩ�13�����	�E��k�ڢ�&i�ⴛ��s`�mho�I�`����c���ِ���(U��hrz�K�hl���n�f�.q�1�Y��0 ���Ui�6�LL��9�� ��{�M�L�����48-%�����nR�r%�El$2X^	cyuUh��m-�hnF{[ҩ(ʥ�V��VKR�1f1��G��%ss��2��� �6|7:�;��9pkfW��#��U�]PR�x���8�&i�|^�^�8�,ܺ���F�2d� �@���I�K�Dc9Ѿ��V�(�uhDM��'�h�f��S���]]VU(E|,����\]]�-�����$'R����[祖Se�Y�ܭ�k2�b�:�^�fq�g�A�"O~�_[Y\�b��M�6������A�
�`+��C�W��T4���f�m6�,LO� �秷�S~orr�*�I��� �3hi�M"]Ɓ�������n��,�b`n~���gq��ҩ<�����>�Q�ܱ����� A"��bA��լHB�uko���_8'HB{[���?Ǟ�� W*���'����旖eO%݋���\V&�%���[aC��㤄�E)��9���ڋtFB޸��1��e����|�8]v��,���Ӹv������� ������~��G���)P��XR�s���q|��C,Y�����O����x����ӏ�J��|�!��/��['����c�|Th�<�|����\�#���G���|�b㣄���̒�F��h4�\�x@���ۏ��V�%=z��o�T��a��Ό�RmN��S�    IDATp`t�n��a�V琎�I(%��B�l���ٗ�xq����a5�A�(�b�+D�ё�����:�<�;��b�j��I��VA�����jF*��T��[�3�X�¢I^l�Z���Z��0�1g#~u�*�?�6�e8�:�� 9͊*�ܬLV	B;뚅��ɢ52.���i-&#�w� 1@ο��'?p�7?�g�����.C�W���ݏ>�������	56����8�g����/��9���`;�x�!t6�q��e�&}����߃�,ί��������%��`����f�8�׀�c	|�'gq}.���Rjz����SX��O��%����8et"^��3o`��E���0�J6Ji/�#��ڬ���l��|*�]_*�7���~[�$���^l^�GĠ�$�f;���5+&�o���M�OL
��C�����4�XD*��Qd@�K+��r�*W�~��l 6K�k����)���rE��V���odĊt�����C�l��U�R����R6���Ħ��p���ag��"�:�b�I������@�!�Q��\��X)�&�J�!�c-�8��D�k�Y�s�Ć����ub�B�@��W���-��V�U��f�py����w�e4dR�E��)�A�(7�Z��b�QNN�X�ӷ:'Wg8�%�M���2�6C%@��Kh�Y�us:��w�����Y�s�)Q6D�߆BU���"t��2�9=�+7&N�����Zk3W��@o{36�7J��W7��3��$�!E;AҢ���6������ylD�H�J�X�"�+?��TN;
����GK�*ނ^��A9E[Y]��{(�$�cޣ��inl'"����L)(������I���<�'��ʖ��6�T�z�,���55H�N�EK�	;-��+��Ԡ8��G���'�q��%,.��������f��alD9����pІ�ǎ�� �[p�+ph%x�:<䱓���"�6������9DY�(�� ����>5�K�:,pZ5i�N�m��c�Ù��3OC�!R=T�u1[�57&RR�YZ�~0�
���߬��co��ۗo�l��y����2:�cK*���
���
vl݌�-�B�`���9�orj�c�KowXa�PC �EJ���ǟ�^Z+r�&#�p����u��ee�Ir��h&���I�;�
�.7z����
����j��1��O�4R��sBis�XX.��Ĕ8ٰ���E{s�>3�$���]eh �.�,l � **T��X�t^�_R���m�����X�D��"Kcf1��5��X��*��7bSo+l�
6|.�|Nq%�,/�e��*y�TB4[@�PBQ����vc��IA��=�ZIZ��zD��'݂�Z�r��:��6� ����'Տ��@)y�O��o��p� ��i��YHmq5��]Ì:eH�ȚK��8����y��_��֖We���P���)��*�Z���o���J
3)�)������ݎ�g�`qv�MV�:���NL����X�>�X@5�Bvc�߅/��a��-R��-f�FV���~ׯ���-a����G� C[zn�;B�=�J����>'��0���d~��y8\n|�����HAx��9|���%7����b��E��`4ABU3H��7�M��pe^R�H�85@a3Ž��)������֓�n���L�:u
�ؽ{������C�&�zx������f��7��������Y+%���Gw#>���ç�+E+�F,.����5�_��w=�(�����%������k_Gs�T�z�Gr���IZ�ִv.��9�417oL���e��A�n��ߍ��s��~�7�����m��3����;�����S6�|l�dDr*Xs@B*��j������:�L��%�qI+.�(�H�-	
Zo�����f����	❤�za,~�Y�/Y)�0Lf
�a�1�Ps��G�+�ք�Q�H�t�z�Ѹ� f�v���%�~ueW�\y��@҂h^@ڠF�؆	�!�)Ww.�v��M߷��/��ǿ�ށ.L���jCP�V���_�ѯ��?�-�yx |��ؽm ��v���w�򮵥�:�{�����5>.�������x��ް����B����V	�
^w���ۀ�72�������$to��F�0�g��YmR��6R���o ��l�X�õs�����B�[JJ;P��7�I�;�2de�%�"�%}AQX@���Ǉ�|?>����S1��1�-�p:��K�e���!���xSK"�C|����SBUU�~�%$�9�I����5'������:u�/\��僦{O(䪀#������F��G��LN�iU�e�E^w�aw9�&�'�����Ɍ�,�-"��"���Ysb,�Pm��M���ŧ���$��
s�G_��i
7�*<P��*^�ɳ�i��`�=�{�|����ani^uN,I��] 29N��Y�"H''�=:)�h�X��u'?�~���+�Z�M�ӕ�������9��� ���1�Ӊf�6���S���Q�M�B46�ZJ��	\��)t*��'�3���8�c���2p�x,�bٙʗd�0s�l���^��7�U;|�f8t�Xyr��܃"h��.47z��K}��6�@��ۂ�~-ȥK�D����1@cS>��f���a�+�v���	�Ss�z})X�~:�K�	�k�.��g��M�2 ��"�̋K�ةga$y��n�B4��������m��z�f	�ǩ	Q���ƀ���ft��ఔ��m�%�T�1�ű�a���W/�����N������j!�q�D���R\t�H*9��
؈ƐHa�t�%A��:v:�Bw�2LV3Lv)����Y��t��6��~�i!�ϥ٨�?��`O'6�ke�v`ۖ>�mBn'I��-�J#�P^It�r�D��D��&eڹu� ZZ�V��*"@7��xO�_K��L�:p��U�<s�}��-ފ�Z1��8�6���W+�Z*���h��pe즈����&�9�GW�nU:�5>bkȂ��rR㤼�u���|	��-~�&�1��nf�H�gb�2.]�� �h6Q�n����n�1��@K�.M$J(��h��i�Ն2��U �7�64	:q�2W���U��U���0׭�F+�2%�"����&�������=�9��~��<��/���|Φ��_r	ja�B�ʬ�TO"����.v�^G��ʽKi��+�I��Ƭ�L*{�!���r�ҰH@��QhʪZ3KC^]Ew�BΝ8�%fq��L"�����7dz�h�5'*r�9���!Ż�ߏ?��Ǳg�4�l��kx��g1qu^��� ������%ҠB�h�(/�oJ�&�oU�Kr���>5uK��V������������^x�~�U����~@h�Z���8N�>K5��i�*֬���sq{҄v�	?���"Q�+_����Ōp$��'N�P�'��7l��\LI b-��>�֨~��P�<u��&���LD�)S�����<�?x�aqv$��<���<��_���O
}���?ڻ�P��J�4�BSs��]�8X�],�6A��:�)s�8���\���\8��%�@A&�+�x�
����c��4������l���VX2I���QI�`6
�z��iQ����`s:�`��*Ӽ�a$�ð��I�[,�]�����c��pf"̄Z�3C9Rcx�ȽSӬ���H�j�yIa^6P.����v�j׋K�Y�ح��XsZ�Ь(5��y�A8w��~t�,�.D�59�#���@�C �5<����V�CZEH��D�����4��WR����3��۟|�W�}����Ԇ���/�����G���lx����A%���~�^~�e8t/�/�Z�����C8r����:>���8x`/�\�N\��"�!���S�T��B��w#m.�g��9�k�x����³1���S��PM6=6�ukZ%;�X]����U��+(&�Q�FᲒs�D��P�X*ʐ���<�Z�`�gϛ�X�b#����>����W�����L:)�}^��d�SS��$3)8��<p�����i׮8p��hm��S=ͮ6^��/��I"$�N.�=xz�z��7����_A<C/p;L� �+���ك��$��pZC��*�U�.Z���!�06q�ষ:��TxH��BF�x���f�wGT��*�Hl}TP���G˯��������e�wy&��	C���~�#�zt�/͋�!���dZ���l��8�:�jx�(?��QRة	�F�*1�|�W\křp	%��LB�k��,E��#�����$�N�����-:$�,��qk�����&�ځlM�:���v�ʉ��$���d��2-H�N5~��7�ڱ3�Z��І�� l˱�*����5:����2�S��Ť�㚬X��b-���r��8������Z�s������3������2�:�X�[ZC"U�f�"�50��.<tIc6JH���wZ��{����A�.6���j�N���"���5Z��{�6����ŉ�0qkmD=��b�(�a1���Ղ�C�z̰kU8��5�
%�aa���z2��/t!�k�Q�b�2	��vw`���|��U1�7w.�]��a���.^C*Y���|�C�6����%�ښŐA �T�Aa:V"I��t]tF�	��UF�eY��\XD4�⾔���f���v�b��W�O/u�r�8��<n��#�t�9�� �/N��g�J�m�0v��u��o-��_�p�W�;"	�.N���q0^���DcK��~{��zBpZIǣ�M-��jC���d�`9�����!(�ȶa�t�%䂩��('�<��D��Ŗ	[�"� �d��������:��)E>��6'�-����j�F��S�cz.M�8��[�`��[�W��B�G�F䋳r�YP�¸JՒ	E��biÂ��(~��Y��SB�"�kG<��|*#bP
L����(��I-E�����۩��uu-�Lj�=;*A��+���=�S}@��U4(5dS�bc����\���x��P��*I����,LcqAHR�z�z�	�';CBk��|"���z[��[p��c��uK���LP6�|=��m��hҩ�F�4h&n�%��C���<�];7IA�.������K�t�������A�B�Z�4��E���@,�y~"����-C�XX����cضm��G,��4Ν����G�C�9	G֑���]��	����Fd�D]H<��<Ɋ0kJ;R�J�@'����k�b���?�m���[�Ù3g���Ol
��ء����v����#��SqU�Ĳ8ya����+�,�&���F	�!;>�����O�K�*N�٠q�|��W���/�#MO��:d����4Ї��n9_#�ƨ �kvuU�33��(4���=�]�����	��}ۆTPX�Yh�b��;՜�[ǳ��>ν�&lv���ž�>��,H�,���V�kt�TP6���n�ƒf*��i�	�s�*��Pցp8)�|��a73�E!�l���Ux��gn757J�������P�Lc>�uQ��>4ː��.5DꙥSfl�������u�_:��z%"ž �N/r�	E6��!����ƺLC�(�L����ZՊtx9}�涿����懶ne��~��7��w~��ߜ<��7?������	�L������,*U�>54|���Ͻ�
~�ӟ��o ����:`�h4��@��7/�"�Uq�c��5Ͽ6�g��� \�M�h.��j"�5�h&����a�
�-pj%d�k���6�o��XF9�]RV9�O��$�A1������	�*	���#������~��x�?$ԆHtU�+�+�qMn*6�WEN8t�8Y����ohp3z{����!�iR@k������z�*�S7.�[��	Wo��V�Z�}�:�����a�f`@��a���ix
p"��d�#�ֆ��Y2�"�1�Nʤ��� Cv�kX��U���PbB1�j�ڒ���f�`61E��,�n�=ʵn�BBm���\�$�L�;�	��)�RA��m��?oȇ��yq��R�S+6C�r�aW]#@!h�iD�_5� 7���nt�..�=}�q��O^nE,B�VS���ؿ}��,ԯ��ۓ�"g��M.���[H��Ȗ����p8N��Jk��b�rqA.��)�:�V��,�;t�n̈^���Ic�t�(22�:؅ݣhkp���d�zd��tyE$9����sW��G��T8'.W��da��ڀ᭛��݌��������#Ҵ���E��=��D�3��^^���F��A*��=�?Z�����l��ldo/!����Yi�x\�̸:���Gޒ:l��35�bM[N����x��uª���T+lv/`�`n)�߾y�q�y�^U���%�h
�9�Ek�)FM>�iQH���n٤!g�JX�D165�����:����o˩M0�AO_+��[����xE���1�f\��Ǎ�Y��6�J�����^�,ત��T�V6��REw;�`��~�����Keu��"�H��qz����vwv`S_v�lŦM~Anx��I����n�3V�~��L̮�br���fq��M�K���c��SvSE��4��UD2e\�1���q��d�1�C��#�M�m��M+éSԭ()�Ë|�
��s�x|k6�T�T�8��ͧ�-$H)'q<WԜD�9�u�2��X��� �it�}Vtu�0�݄�'�L�� ��� ������WQ�Hϳ�����uN�+j�t�K	.���L'�X_[����իrX\0Q�dxI�-��]R\��iy�u����x�����S�kw���<���sJ�P[�����ӄ��2���dH�eKڐ8�V�acCD�j�(��",#�D��s����籶�,A�Z�7�X:���`/�
#�Sʦ��XŽ;����ǱwǠ���*Kf����-�9�p�o���U����+�`=+��cJw�{8�}�"v�L&��E��}����j�#W����S����+��^J��͉q�U�}7Cػw�8��!�Â��<��ዛ7o�fu=��%�hmi���{�3��$���-���+�XZZ��褱��`":�]%�K�
Ai��aF<c������K��P�#G�U6/aoA��~�>|�=�JK`nՙb�}�M�p���/�ɤf�1�~at���۔�B�YDFI�(�^Y���1�=+�����:"�7���Q�un
�2���,�<z'^}-&�1�C�!��ad�W�%�4�R9��0�*�v�;G���q:p.��$���5��wa�.�-�&����_�Bf.�y�(>�0Ѳ���h/>q��3(�ƺP}!��94�N� ��N�l
�J�Jۜ�x�(��з���^��N㯿�,T-��	���b�!3�_��܂�*���(3��(
�;�XK<�}�k{��?���T0/Կ|��ϼ��[�}�=�>����o��B��X�N/�P�2t�˹"�]����Y,���hᔵ��x��{�}����]g �ZLy�����~�L��]�~~I# �o&��t�H�ݟJ���&b���"M(��[{�$���d7�r�%�t��bwH�oHRi�'��ȌT6#c0��N�߳S�z�7�7�ӟ�#Y�J���]����!�"�y����Y� ��c�֌؋�#G$�X�.���ŀ_\h�,�8x��-�M���*����������~�#o���� C�d�c`h'��� ��V\�YD�bÖ�[~�sO2�P|Hzh�('#���$��Y���X�Y��U mHd�=Ey�+ꄺiH��� =���&`*#BM0��N��VT�"�
���HC�kJCMf����*�>I>e�B-m��3����ԂZۄ�ɪ�2�ޔ�P8���-�72i ��6S	[�[q`�ft6�`)P��.�M�f;9`baק���!���I�
��a�]    IDAT��T��V�asW�ݹ=�~8,��P�U��F��D����~�"�x�,���ymZM�X4\�>ԃ��F�\R��U}���M"m�쥛8r��oV75��"7�\�B�T���GGk=]����PpL_q�G01$�c6\����I����e/s�X��`GH��}�pjE���8��3�C�	���Åp2�sWn���+(t�hE�i��k$E<�Ex�:6�����d�Y���'��O����o����f�.���h�J[6�`��t6pZ`3�-̡��!��	��7�p��,G�0����f�o{ؗJ�)L���D__+�6w"�g�H�y�{ND�E�q�*�ߜ����铜	>���c&�1�$��"��PF�������F�v�;E�+�sGa�I�I�pkn��]����\�>�vwb��0Z�9���!}��	���=�T�6��.(nD%#���-�س}P]���S ^4�-�qe|�/�@4U�ߓi15`�:�B�æ�f�6���V��t	t:�'���.�ss+z���Me�](�����\�J�M-3�]��� �` �C,E+�,R�vܿg+�t ��D�*|$"4\�9���X�,�޹��M����̴��2i�!@B��&�������'N3�lFʐU�b�̉��T�=��s��u��kR�	�7	����,����瓺�s]? �TC!u�H6)C,`i��d_��`��4���[���n�����
�(�n�43�Ks�����t��aҋ��:hl$"��uu	b�]�#�4���>��Ǳ�ͽ��XY������k�%w4����(�|w ��p�Z_GE2��B���l�166&nDx��ڜ��Zd�9����oavv{���'?�ii:�9��G� �}��8~���d��G�8{�,�9"ַO?�����u��-�G_��/S6R##[�/}	{v�������`�B,vAPD[�3]�z<�!g���M���e���I�ꕣ0Ln��S*�F��ؿ�w�v	x�s�5�;��;�C�yU��M��ep��G�Z�&�T��ƺ���0�iBt��@j�8í�#�IciyS�3X]\��
t����^�$�@ �P���l��/��/ ���[o_A��@�MGvi�D��*��)8,(�6W�eh3�Hm��eC {��J*+��DT�$D �t�b6��*A���X�d��At�Tr
���h�L���ᦲQ'�tPi\�w����b�� CB���C��� E�a�`��%��kJ��D�i����������G�.�ח�a"��a���o�j�j��P��z�x�m����
Y�8lK����������;���^y�Ͻ�#��i}�����@UDO8�������Jt	�?=�=LN�I���WՄw�����B1��,v[<Q�[%�8m���o.�'ϟA�������r�!੪7V���@�*,�$�Ƥ!H,N���
E|�:�EĂ�BH]��5	�X,�JC��7�Ê�e����;�=��l�y�U�-�����Qn�L6[����ĲkeiY<99�{Gww��&����^:O��)����.'>����F��������?�`�Q�Q5���ҋ�{D[�0�֢H����`T��	*I�������"b9�UG6����,6QN��Dڕ��}���7k�I�4+3C2����Ȇ@6!aQ���0/|ޥq31�&>���	�{G�?����L��#S��gY�&vѴ�#�Qi ���
����!���OP����:�~Gl��'�v��Uib��T���ׂ�;�r+��T3IfXuˑ������e���,��(�ch��,g1�݄������Z��.if̯$p��$N_��7B��/ݜ��bd��Ў�z��H����X\M���k8ui��_�LXY��Mr)A�3�~6��a�� B�TT�A���͋\фT8v��\�@��{T���!Hn���cþ��ؿ}nk	f#���%b9���AD��
�l��z'߾*(����ۈ�A'$L�&�g�V��lK��U�e_iG�lťks8}aL�74Zh9k���Fk���?�[�t� �A�P�*��`�9���i�tE���v8m>h�B�؅3K��x"����`P������%ߟ��B8a�ͳqkv��$,E<�q��C�/��䓲�*���2�m7a��#[���Hqj���,Xل�-��(���1�=��4]�&C��ؾ} ��_���
"fs�l����I���S��i�ɰ�
\��:��D�ژ�C��};EoU-ӫ��V�:�����g� _քf��xUs�I	:�Fb�H���{l2�+�2>'֥�d�\��زeɍ���D�.�E�[����	��\�9����X<�$�+0U3�=҇w�݆޶�&�n�))�9�+TNqi|�/�#B�*��/$Ǘ�"6p\ɹ�^U��V��*v�|�B��ͽ������R/��ڑ�'�u���̀4Luה'X��6��hV�������8eV����I����&�m��;��@B��ѱr(�@:ZB��	�Y� ��:t�&ǁ7�$�|�&��Ne���"�)>�N�	��[hphx���}�~�B�
����̹sغy#[E�����ZO&���A�b�(��:��ɤ�D2���E�vب|�������-�-�СC"^���z��/_����Ͽ����K���O}�����mH!Oz��=��^ý��+T$~0����C��(��<v�w������p`�>����,aiaQ��Ĥ�FG�j�Rr­���c�'&�L���D8|�"~���Z�(Rɸ���z����x���R��,��h/�r'N�D{{��Al߶��ZH�L�����+/��+b&1�u��މ��.�|�80���\�(��ff�<?�D8,�y6S��5����l�"��N��yud�x�b7n��ϣ��L�W�r�p����@�sq����Nd7��X#��*�9[D9EK�b�"�,C"~��1���B�j����=�t5݂��F���+{(k�P���Z���Er[�Z�^g�V䰎�*
�H��GQN�H�1�V6�;^٪#F�]g#\���e�Ø1l����א��Prd:H��4p4�͢���U%��(g���&���������o?��C���|��S���W������ں[w�܎���V�+�.�"�&�_�W3.ܸ��(�M���x��*��;:�v���n��+��� @��q�ˇdՄ�^�/_~�f['4�/�q	���yr����f� �2A�
H�Mcy�f�/#�>0w���k�4�Z��+�N&u�7K����2����ۆ���"Vzss��YܽwC�9>.�Ȏ�jqJ%���♓�NkO�|�af���Id��W.����*���$� �{{��jD'#��Qc�,I�V8�>���x�����ah>�B�:��bp���E$�E�q��Қ��4-��������s���H`zl�E%�Sr��8u�Ee�l�9�.�S�$.\8�a�ؔ�J�'�eH����U�ze�?������������'f��F�H�������zC@�`�!P�r�7 bz�����SmڂJ�8���L	�IY��<k5���f��Ak�	�]q��U���qƁ��"��uc��Q��ՃB����#ڠD�vs�;!h�Q �O[�n���"N�����e�,*E������h����t��	g��i6?E:�)
�ba%�k7�pki��]�,6�意��9�Lw���ɋ{vmFw�F.�Y�>X��r±"�^���c���F�@��T� ��c.c�`7��=
�����߭����Y�������q-�����6>�B�b�h,=���f�¯��j���1`C�G�/Is�����.�M���fA�\��e�H��	ފ�6l�*\6M<�I�sy��Z�k�Q�v�,��@�:�����6C/^e��G!Eow�nߊ��6iN� 3P���+�Y
�l�
B��Mx��AP��P�W~M�qR�.D�8�M�VŦ�fܻwTِ�+��� 1���0�&�'�t�O��AI ��@��-C����ǜ�����Ya�=(�-�X�o�<�\�.�G3a��f�aTs�x�`�A$c��u��@%3��p��k0@6;|^/��ҋt9��}��6���� �0���x��+8uaL�S���3\.7Z[PHe}Ld�(W
��jǁ�{���*V��Dc7�q�Ҹ؏����f���)�hp���waǖ^UT��Z���X�&������^����O�	&���F��Ų#�H��9%��p�Ά��hXf�e��Ÿ#���u���~���������X-��6�o�"(�*��մ
��c�sU%�������� /�|��2�b�*T��2O"�t�
,:���0rYh�B��=.�N�:>�m�z�d�\���!KAj*)ÜL6/\{� ��G�����'��][�� V��Ϝ�񓧱{�N�O�%{���C��������%`n~^����ߝ[\M�Sx{v푠���*^=�~����^��҄O��"�}�7���](*�'_�{y/���]���{���p��a)�yNZZZ��3�H�ꍛc�ɏ�����@�ğ�����\lɗ�ŝ�C����^�|Hvy��pe�Ia1�u�c%U�/��sGN��n4���4�~~������dkkzyϽ��_|����#=���EK63�X�f�����_;�x2�` ��"z��4(Z���.�+�lf16a�a,�*s �*՜)�C��P��-hkhA��D5�-��¹K�?�64�1e3p2�/����5���m�1e�E>G2�!�&ASY�2J�F���\����&����MS�T��5 S-��󠥳]���I��ӝ�3��"m8�����F������K�_��h+O&Y3���ќ"��6�� ��Mh��\#������C�c.�C�f|��#���Ͱ�^����z+�(�'"��#}��<�s����������[y�����P-gd�a1IN`WV����u/Vc	l$�By��r�����ڌ��Vl��@�Gx� ��<:MM�.D���ǯ��×-x`�Z`��n7u"E�\��p8Lh�2:���4s��0�@1��6�)�����+n�lv�ȝ�E}.�,悒J���P?z���Z��;/0#�ޞ�nI���?�p��1
)ٵ��b���Q��oD��������v�g'Z�1>~���hnlAg�KP&�����ݺK|����boC4Y~�"���3���M�ҹ�	u`������/�W$�C"[^9E��Q�]�Զ��	���#��:���"�ڀY6��N_,�*
ʍ�*n�/�(P|�ȁB1��QB^�ǩ�g�J�A
�Y曤!�ǘݻ��?�1�MN���)��(��@ؿ�-�C�������Vx񦾫ؿ3ySڎ�F}��,4 ѕ �ii8�e�ta� ��:\�?
��C���p����c�Hӝ���@:�,�D�~��x�v��Bw�_�	�)S'@��d����8{�nN����%lx�{FH�q��g6�%>�t�0'|j3+XK�!�&)�:�&sfW�nF���l��;7���MTH�To�@��N����_����h�0��
i�����Q��8��8ԐZ@��4ҙ�����d����(�ܘ��F.o�Ь≬y��P�z;[��ф�&7B~�Ej_�(V$R._����*L](L����;z�w�_lFy�r��c�N��X�څ��+�̕�876�X�+��ph� �A�B��f�qD7��Æc��<���*XZ�ҍI�-GP2�k��$�3]��ǸY9��T�4LP.�n�(�����[�r�JȺ�&T��Ao�ML^}�$�\��!�|o;08�*Bۀ���DFYZ�z-�.���061�������Q��yp��z��e
�"�4��|��Wq��5�"���ɱ�Ԅo[���^�����̈́â�KJ,a`f1����t�r�Q�`�Iʳ��ߌR5�|)����7�2�@-p��,ο}�\Y�W
�=l*E������v��]Є�S��jE&���Z4����qL.D��Z�\`�]�Ю��2��u��u7Q�KZ)����,��07/�_���wB��k��:�>�]m�����j�=�?Y�׬!�+���k�sR�b���"�BQR_h�-�i��fhMM�4H��Ƃ�(��k?�̭[2�ټe�;�TC�@8��D2)	�d�`���k0e6���_������B���ͷN�C�%,�]>���NY���F����c�H�0O� KKXXZT��\��By���'���m[}]X�ǡC��g?��؀S��/��q��|����l*�/|�x��GI�x�"�z�)l�:�cǎ�'?�	旄����~����������}\�zEb<�_����SO
�oea3���K�h	�j����2}Pī������P�F
������//�����i���!ې��j�����+��|�*���Q�^���Çq��u<���xp�A����hV��Jd�t'�>��gO��VW[;��~��n��0��bA����^���Z.#�-�4���0Hŧ�B�z�
�V],���
bӷ�~�&2��@4�B,*5���,��̡��	���SG1�B1�����gOf��RJN�"u��6�-(q�v鰺ݪ�-�%�(�ϣ������`��*�;���T�΁^� �~&�Bv���-�%��	ape�1�8AQ�@�"�[����-u	�ي�݊�߁|S��܇����t���|'.Oa&�D���@�6�f��q/`��Z�z��֪�Lt5�{�������_���!�Y������_9����U���+�Ų���ӁͰ0��N �wMfX\.YD)��koŖ�NV4:ut41|�S)�!�6Q���&�x��4�,Eo���H\+�F�B�S}FE�\Z�:*��\=���K����iX�?��;H��<|���u���y0�  "$� �"%K�hR�,˫��v�۽��=W���Y�뵵�h˲�`�E*�""g�`0���t��u���릱�������TM0��~��}�'��ȣR�A�3��(�	v����hvg��g�͂P��-ؽs;���#�3��%��k?����R�wtw���IFG�p9=F1�dׯ��������]2�(0��Ԇz���KF�!��\>	�al6ń��6S��1E���\�1�^�Ŀ��nN�J��B�l�Н��o�І���e1���@ʩ�`!Yg"9�HK㳈�,�M(�,lւl��bZ,�ذ����"�����H�[���	��)��a�+�˴٪I	(��Q	.$�؉g>�	��L�͊� hn
9�sL5DB}�T9�5��*e��x�[���M�Ws�m����� ȆM�OI��R��]=80H��Š�#'��1����y�N��$F���E�����L[���ף�����d�%~V�ŉD���\���RT�|��9�Un*��΃�;���݀��
��.�<p�&e9*&3�bx��U�.���T�<A+QҗY�F��sP�� ���j�bW_;�������	�l�ye֤[��m�xc�F'��X��X8�e�M[���6�-�źU��wy.�a�!D���6d�e$s�.m`=���S��f���<"�1�)���7d�B��ҼpaOf*�g0=��D�(��N�(=/Ԡ}�]����d=�6��[.j�d+�{1���Z�'Ocv-w]=T�"#�Y̛a5٥����}AB�,z^�ʇ��Ag{���ͯ�blj�k[����d�ߧ��cⶤjV�dEpωYɘ$����04�Mr	H-c��+L��iiZŊ�p
o�wK�Q��A0��8��������+"j6��eJ�X��F����)����P=A��I�v:�2h�p��~tw6�ZO�1���u�h�h��x�<�X� 3��Ϡ�k��n���    IDATFo���y��ͬ�)Hg-،�p����g�q�_x�tL��!��/#WLK�4�ͻ�;ѳmb�Μ���#���
��Rʕ��!���>�u�_�\I4KrV�" �9����u�F�(1���B�@�(��YK��y)�48������Y(D���1�ŵ��3��*^&���I��%6�����Iem�@���	����j���I�q��~�@�yH C@��&Re��� ?�K�IM%�r��uY{͜>�����5.�U�Fg�CJ&�D,,{Q�����4����4���2��Sh�a�[��`#]2á���o~���da��wN�����4Yy�CطsP�`iTĞ6#�ߠs$��O�D�ˆ��x<G"�#�&���ԇ���FN���ʞ���$�ߗ��e|�S���s���ߐ�ɧ^�$�����01>)+�����?{]�}�3��}��'��_|Q�ǆC`�������Z�Al��anj�tn��
\��U�B�u'4��}�I��:�k���-|��7�ʻ��U|��=Bq)�#���x����ǿ��&�y�=N�E��[�`qs�}�q��oC*
��-H�3:v�lE��Ib��Ǐ���6������2��0�u��Տ���B�L�;-���MFERA\
n[>5����O���%����G(]M��i���/B|���S(�ҰS�+����1��#��Ƥ�"3`x�p���
�B��SN���<�Z���i��. x	���dz2���ӊ\k�����z"-Bs�i�hh7M���j���d:-�i���
{���Of�V3N+�~�w��{aھ�^�+���scSȚ�0��`Ai��9݂����1�&��+��d8qx��������7M,�����_LMy���~�'g�f����2;;r�xA��'=c8���L8;^�1(���M(d�ho����@g;���p��\�]eqB�P�ۦb3U�{Wf��Ϯ`=e�2$(�I7�E܄�|r��58�
vq�>���k�GWyd�r���md��J�����OA0ř����s����g�N�u�a:<�Ӂt!�w���p%7�<5��ͭhhh��9�!�&+���Ȩ�ɻ<p`v���u���~��u?�ۘ�	��hٜxs����.F>��&��8�����x����k�`u3]���Ѕ�w܋m�ara�[q��n�T7lVC�hT�eTL%��t(&�	��-"�� D7a.�a�`V�(��m��+5�7Gx��*D�l����.��&S3�e
L�})�Y
�K(�!PM��?��?��43���f��@�>���E�l4V�����r��!�I1x���@���Do������IFIC&�����.��68�eT�� ;&�ɌQ�_���FEFN��ڄ�E���MA9�CGOk �-q,� �ת�P��`~-�K��1�F�bL�<.�k�6�1�ӌ�z'T+}�F�bw��eF�Q�-�\���\�V<�'��e��|At+���0�TF�931��,zZ���ӌ����i%�Hg��h(����V\���Vb)XL6���N�TH����߆F�CB�h-���5C*'y �o]Tt���D%�)"_�be=�KWF���	��'E&|�wbGOTGE삉�Db,�ű��o}6ʺ���)/Ͻ��G�v�(Y/��	�R��ݴ����W'��{�,�li�ٮ�� Q|�����.�4�[�L�#���*�6G��bh�\�c��>6��p6�q�ղ.��GWD�De��6q"�d��K��#��b��.��э�05�w��Ya����;?"�|��/�L:��5���h�[נ�H�U%���	[���Q�:%���#�1%Z�V
�m���{��+2���Y���k�@8Uƻ��F$��D�
���	��x�����"V�D���&�6$����UI�.Z��)QDS	�S�UL
KJ ^�L����f8��Wo@��$��au��IJC����[	��5��C;Q�J��$	�*���L�8<)ӮH��;��'�v��(UOr6����H���,E"A.�bE)��b�(E�L`oK�Mk��6���O)���S�k4��:���"�m-Ь���A��E0ς�v��S	)��Dt����l.W}βP0e��ײ4c�r�z|��o�KNk����361)_�z�ۤQb�'v�EL&
[>���z��gǑ�;�2��5�w���7�m�x�cOc��>��6;�I�ϭh�j��}�	�QD#�x܃A�� ��!�����w��7�|�hT�r_��o᳟���}��!-�/|w����2�eZ@0���o
���=��G�����6,<nԲ<��x�ÿ��ۍ�Ʀd6�8C�����0-�5x�&3Lv;��y|�>���E�Ã�s���+o��gG+��;Ĳ��CE�?u?���|
LF����ޭ�u���/1M�؉�j���1\8wׯ_���
t����&?q��P��-��ԣ���Q��'�b��A��8>����ni�$u��2W��L��STR9�Z���ΟG|j�H^���&�#�si|�_;�����DL�ي"	�G�I��=ё����(n��nCA]s#lM�@�G�ILR�ayz�Dݻw�]w���H�T40?�u6]��7]\AauӸoB8�~�L�.ag#T( ��Axj��!�a���bE�$m��������q��a2���8�w��D�k�
L%6����,�4jM@VS9K9;q���}�����3zc���>��������k��ڭ��s&#L"<2Rj��hV��kb�S��e��+�B�iV��{��]���"�d�4��P��3O\,�KC@Q�J�\�.�J|�瞣?jXܠ��ݮ�(2^����X�E97�q�&D�Q"�Œ��E�iw��eK,�uSs=:;�q���9~��R,������6<,����/X���x}��/���a�Ӷf�@d�TBsK#�]��p8,�Gc �fxS��8qP�V��r��(����$�D��?N�ngQ��/�|�EL̮CKW`u`����8���D�X�^+%	�2�2��.�TԄ۷������ڄ���՜�4���pť�b2&��B<�Y�#mM�R��Rj\����V)ƈ��BX��OXw��94��~��"T�Y���7q�TA��6%��?G�^uBPv�m��[�G-3��{�i��jn�R��J�T�bC@W��EcЉcw	���x�NjTΠ�8\�5>��K�S،��p.�6i�XPZl`9������Q���&�{m�U�].�KV�,*6"Y\�v7&�Y1!�q�5��z�7���
Ķ��p"W2c=��������� �fw�6'�n�l8!�n&%gt�Gw�{�ڤ����I����q��ȕ�ι��^��Z4��#��IF�2���A��7ë*0SP8=bG�U������v"ON<��y��ztbW��a}#
�נ�1Hl�`���)2�瓈���XX� �,��pI�Ŧ�뵉�ضF�꼒�@���~�t�ҭp���s�����$���
��p
����P]���h���(B� �Pȥ�K'd��mk���>٠nN�!�Z��jL�#8J(p�a2�G:{0��G��1U��v�w�;���3�&v�V�-.9��\���،�k��3Y�)o�p��B��t�H97�\M�*6+N_�z8.�L��N E��m�Ю>(
�FUI.V0���释�oL!���,��2J�,"�kh	9��Ç%�^&�"T�
�hFV�!�S���a�35�J�U�Jp;=�d9	*d��:�:���)v�`3���F��G�9��x�f*IC��َ� ؁���!,&xU����
.^����"re��q/���6�wp�fQD�ς/OJ��� ��[6R|��J��9�q�k�@MOR+�k~�RēҐ�!Y��y;��Fz�~V�Ԛ�?e-�m!����42��������ȟ�^4�G��ݧ��)`��̣M���WJ����'�fjnN�I���F3@*�b��!_{J���R81ԏ��q�&z>���7�g�����x쑇�P�C" �Ev�X� N�y�T�[&��C�_��1t�h�;֖�F<��#��c�1��w�F܂�<��}�w�>�����w����ٟ	�ǩ�=w�-����M|���{�w��������g�CGG^}��x���f�l��!b\N��^����A[Sr�	yR;�
E%��D���Ť���M흀�8��0���|��}mF�=b̑�/��ц��_���`a�h�{����K�������4tt�s,�Έ~� '�%-��w��/<��m=bLJ%�2�$��<�>;�ӗ�bzn��*v�u�3�x�;��ہ��5a5�Û���lhFС�Ò�!7?���'��[��PD��/�!���x�9�!}�a�'�'�E1�Fbe�Ur1\�&"&���}���ɤ��g�W��duM�`
�,�+(3G&Bѯ"NѲ8*��U8�d`�P=N�8]��y�:�Qt�� ;z>>ǢQ�@K6ln ���ld�\�dvN7��X,"C`�����:ǞX3���o]���	�狈��H�,J��,2�L��X�MF�!vߑ������������xC�_��㯝���͒+h���B7��I� A�[s���y��h�CA�B�*�&c�p���+�}-�mnB@��-T�nhm�310۝�$9�Z�_~�M\]G}�^iXd�a�,�bf(��2 ա���qi��3�RaiH���cwR,��p�l�;$ʼ��}�{����N%173�υ|�1<�����h��x��ױ�4��LNR��:����'�}�$F�]7�jZZea�C�D���8r����+H$�%vh����֌v�j�J�G�� 2!�Ƀ�LL�b+�BCk7z��`x"��������d�
���������+�|�depGg�۫��P�v�b���G�H��c��(]�͜A�EY�П i
��9 ;Om�œ@��,l%%��!ŖUX�V�
��CAC��3�;���~R�
זl:�h%ES���!�P���ZLP���x-�M(���>ݒ�I��*G��)����7^�%�f��p��9�-A:�~�'��I0��)|�h�dV�f�]Լ~��wc�8l%�u5�Cy�u~/�Ad�r����0��%���U����qذ��	C=�k�	'T�d��
(3}Ru!�W�����z���0��%V�F��r���H��11�@ո�J�,TKQ\�����~�Y��"x*(ea��qitF��k:MyP�g`�q���m��S�\��qv J�Z��'S c�E޵V6����VãS����# �0�w�]ی�R+eE���ƍ�3X^Kʤ�E���@c��]M����"���Q,��v���J�υ뷰��@*_���X�ՎR��1��`�i�¤XѨdPP�VB!��C1�Zĉh�X@���-vn��0k���RPh�&Tҙ�%3K(Ilko�m�uh�M�d����c��ZK[��ES9��.�����R�����ط�]��x���OB�����02���~yZ,~��z#m�jE��Į�64s���n� ���o6�ܚƹ+7���%N\�2�R�lm�!��ɇah�Kh�i#D�+t�p`t<��SX�$��	ba�ˉ>��NhI��xU�dsi)����&�Z�2ĬR*IR+�%�R��e�1�Y'>��!�49�(
5)lDs�^���s��ȗ�~Eq��i|-F;�/U֙�͈���N����o��C���TA��zJG����$���6<L�Th���NI�%F&#��n$��d���g���!Z�C��D�H�%������F�A[�~Wg�4460!�ڀP�$�F�T���&R�8Mgc,��ٴ����u��Hr��m��報7��������mB��x����3O���.��>{����	�N�B/�05=-��������:���EP,��퉈t� V�,�:ۛ���`�;T���ɛ���'���՗�(�⟽���/�B�Q��=����ocjbR4N�%t!���@Pd���cڃ���x�I'z��'pǞ=h�0;6��[c����X&-�A�I�45�d�����咯�P�� �n,n�/�~~a	�YC.�{L�$��|�G��c�¥�������?��WǱ��
5�H�&"PF��z1�;�8�/񷰧ǏD
����܂L�n��av3��H\�Xˢ�͏}��I�_<{
��⧈����܀{��CwE�b������k�9��5x���f��`�b��`^��N���4f�#��'�ͅ�H-@���AG1��l|�3�k��H��3O!�P��hW��̈́�^FN�_JQ���E�Mg;��G�68N�;{$�SDK[]�ׇt
��u�Ӏ�df�j?�u�8qw����@��q$<!�v�~z�
V�D4`#�GI�Ca�,M"H��2���+91H������+��o���]C���ɟ��{�h4��^�d���ĉ"W��33EX��RB!O���8�7�����@>�Svm�Ů�^�Ȑ�2� ��W���ؼ�o��[�xsCrt�[Dŵ"���T)����~Cp��[Hl�@c�V�!0��y�fp1Ul�	�⤣
�H��.�s�������������E]�!����~�㗑/dQ�� � [�L&+:���� /^��q�˩��$�D")j��:
:556�$�\D�P�F�����a���p��ゴ2����+8{�2|�-8������~�?��I�*��!4u�F��!�6��dSy�ilPU��BI���,�|Nڅ�N�a��5諳0�(<��R�eZ]�9��	�n R" #�dc����!/Q�Vl�*BN]�FǣA�����q�~<���pxT�//�S��4��X�0ʼ����J�������FvSx�O��ڄ����6���j�_���0L��.�CCh��a�+'+eC�N'f[�,��N`|v	�D6;��jp�D�g`5�"�mo����E�=��$E`p&E�JD���-�u������ց�V�DRR�1�6�ْ��2F'Wp��-$��m�$�0d\���MJ�i�vŠ>���f�{�۰��u.��w�`�� �T�y��<:���MY�d�@��ӊw�G{��� ��Py�S��/uA��Y!�ɰ8��l:�a+����
&g���{+�	R���9�F���jL�UK19�&������~�6���8Iᰉ����F:����qA�9f�6�K�$D�D'�Rt͒]u���~�,f�0� #%��mX-yL)��� uI�U3/�1���� �ƥ�%<Q��s���Q���`/��;Q�"G?)c<����h�	��v�dAha�6�F�s[����+$��R.�hd�dn��&q�9}�"�����C�PE�IZ
�ʒ�A�QU�������[�E!��FѸI6�|&�T2��?=�{�;��r�K7:R�ؔY1<��#Xڊ��&�j3�>x��I�Dx�������WdB��Qp�h�������ht-�������}t^��|Foj���ln�ob�֢�E����4U�Y��p!�ÄH8���MYc$���Ⓣ��S�3g)����r&�e@V���fQ��jr)�ǀ��'����}zdբ�F�	��܁��i��sJ$b���]]�g� 1A׋�x�Ō���ګS5r�(��')w��l��Kpi{�PT��ۼN$c��1,̪�����p����w⷟}w���A��/�Ͼ�q�;z�iF��193-4@������rQ��ghV�g�F�]55��}x�>:| �s�sb�������2Ƽ�'>�A���[��׾&������3�<#�13��k��8{����@�������^��$0��b��婧���}�r��~�n\���;U�8��ѭ&/TJ^?.�_�-��li��Ҏ��A�\K�ş��k�F�ѽ"*�DE���N�G=���q�hP%z,r    IDAT24צ��~�_�A���[Z�R/H[�lZ4!��]��>���{��ZJ����*�����5�.� 7a5�q��a|������k��#�L����G������@iq��X����&�`7)��6����V'�ȲPQL��x�"KKp�e��U,�ZIsn���[�p�S�fmWd����T�U+�P]n�%?�kr��V�,�Cm=����+E�2ӂ�����V�Kt�bj2Y�:<�~�S!/4:�7m��=b�bF�jA��B���h��!��o^��߿}7W�X����
3�Bk�@��؂�L5`J)�k��?���o~��W��h���~��^�Y�o�a��nǪ����U���Aie���F��,S��Fس���y���|�E���{���S6���̴cs��ZQ� ��Ƥ!�XοLƆ@lF͆�Q~A;M��ç�2!~��FC�	�� *tE��&�"M�tv�-�y���u�c+���c[o>��s�����5R���<^��Kk��܌B����M� ��y��{�ލ)�@�͆����X��'�w�^�n߸���7���K&���;��C�J�7�d,.�����d�r`p�1�r&��7q��,2,p��Zйc�,"���4�Q�l�+(������еfFưx���I(H�(P��bJ��e�O4���1�j�,�! �KA�b�b��2�Iڬ.�&� �n��8<b��9����T<�8�Lΰ4+��0J��,��o�2�O�	T�kH����ͷF�}Bp;��Y�|�Z���� �{w��=�������bC�d�����5�<ܞ����D����q��΍�ۊ�/z�\L�$=�h�re#��.�`|a.wP�h�Ә����u4��EL�~NY�L�r
.^���Ü��n�5(�m.�Ɔ@��P�x5W�E6v���ی��-2!h��ol2EH�4d�fl$��82���E�+�1"��9��]���%���av
�I�O����)wc���G���6;Q�Z�d��f�W0��%����{qh�Nt���Gg,���-��<��eR�hu�#T������kAO��&D��<��#cڕ-��\����'To6�[
%e�H
#���p95��mYoH� U��7�S|JN��J*+(�	�&���b#ː=&AKfVɠ���x�+�rPIÆ�4�݇z��J!c���]�;�q	����6�Q��`h�=���N�S�)�L����)�����[Z��i�A�>�BW[�dU��Y�f<���9ܚZ��V���U:�)EG������2�y螽��q:��`�m����Z�ijE�1�0QdN;\�5��@Wo�H�����8u����L�t�]����d�����3�"�֠����ݒM�����Q:_"S�T�+�T�`�q	:bآ�1��q�ɔ��t�!��t6RE�5!�^�Hv���-bm����$��j}���=��Z��f�?'������&0�ю��f7rj��l&%nr$�B��tZ>'�*�#�6���p�D+F��JYl�Im%}���F��	�)�Y#�xF�a1kx����ۿ���蒢2�/���+��������	�ǭ"��a=�eP�vI>&��|'^��H�tR�_"�}��@��z:q���{�	i~H?b�ط��[�'@�.��=��[�я~$I��|�s���� L��/�Ka<���x�t�N�>��#,`��<�����'����{�5+�~�.�:�R*��.�?K�";�I1��0�d�b���jES�LG�����s��*~8\~b�<��%|�ރ��'���:5M1�����^��g�#I����baZ��QD[��a����to�#됉��lN��� Y�T�t��A��1�Me\<w�t^����8<ЇG�A��Bdl��א��B%��5_�E�L�"�o�(}�І������H �����:z	n��QO���)Ф� �Dv�|Fv��W�
�WF�,�$UZ\��Y��
�M!��4H! Y"��ʀ49^uD�-
�ZIN+ٜ�f�r��Ow@���F�����`udt ��P���{��?t������?����Zi�,����D�d�1����*���=ۿ��?����Z5�?}��O���}j#��S�~Rmk���wɫ;+��E������ؘ(I1�E��{3S2Y�������X]�ՋQ����Νh��!"���
��ٌ7ޛ����$63*��>I*�!Q�+[�Y�O��knHC^��ȩ@|m��&�%�JJh ��2T���v�ai�G�.�Ć@�;R�ޱ�}�Y�n,�$��q��i�rC�f
2�'��ر��o�.�ꓓS�F⨫ɢǋ{hh�9�Â3g�㭷ޒ�Y��@K�O~�1l�ކ����el�#�/�[���&f��`pl$Q��̊�UO�:Ѿ}�d��M�&���+��UQ����]n�@,MLcs�ʛs0��E���H�uf�P|��ʎ,��"��11��V�6;�,F+f�L.Xl�?���p$��b	�RF�ѽ��ouM��]��*��y��1���%�¾TE�D�i����ܔ	��q�B�@&�(XUGp;�6t���^�qw[��wnÎ�:qB>c؏�aF0��)Mh��$ʠ�G�R����t�l��Hl��s�(x.��ؠ8�،��Oadr._ N�!�����h���4�-�)9(&M����9݅�x'���Ց)�s,
\$�R޿�w$��I�1��,���N`����w���A))*f�M���p��(��Z@��-
4UD�zd� ����
���czfN�A���G�]�]�*5D��d�Ε������6Sb��
�����v���MA���e\�X|���lp5�׹�s�{�;�2�TH�*�5���d�o��
C�&0�E��YQ*[��#ݑy,�t8�v)��|I�Ȧ2�ςR.'�i�U� &�,�����LDpǩ@��S
Aխ�u'97bJŝ� -�^L���mx�{P�t��e����U�.�g*�5+���T_:ښ$�E%��
f�y�%	�7��fq�ʰX��h���C�l�#�	���r`bnU�	+a�ͤY���)�$D�����u���C�򋑩���E(��q>֕�Jf$��0� e��J����n�DGG��-.o��L�.	N���$��,~��^���~1��� �D_gr�8L���ְL7e��KNx=��&�K�Ҷ$��[�Aw��.�x,)�)Z/�YF�/~YX�}M�*�RP�*M���p��T���W&�"�7����5����j� A����W?k���.�����Z+��K�}S�8��J���bX!Z�����pɒ&��M��
��'��Ϧ���L`��!Ј!/4Ҍ��z�����'�o=���!�O���3��᏾�Uq�ڽKlf���Pf�MI�T&+��Ԕ�X�)����#H�b�A� �*��u��=��C�eO%����/~�Ν����@��P��̌L>X�?t����a����N�<)�|����񜛛Õ+Wd�g0'�c��ă>�m]]p��ũI\<{+�3�|�I��n���Zb���M��ƚ���P<�}��������cЬ>X])賙-4�<����3O�M����f�������1~��I	6��]���~k�Z��V�e�%�Km���9�4��w�h����<�bZ(�A��{�BS}�Ъ�+�Cuh��ޢ��ㄿ\Ajv
�W�YX��"c]��j�@X9��"����]�>�E�VP�
C��O���&Db�e:D-!u>r��_�^��PrX��aR8�9��A����5��c7�"�4�P��~ev�jC�\@<���#Ќ��2��*�.�:\^����������.i��hn���~ J� �M��{o����ͪJ�&i��f�$�J�!�Y��������_�̯������m��Ͽ���x��/���qܱ�7.������azj&�P|�(}&�Γ�5�R���W��X>��G0?7���a�>ڳ�u��:U�|%h���*�<5���"�� `iEYq
�^K*�PkT�	^8-�4��N#�<�l�	��"o�QA>�p`m6��t�u������)<��	<�����B$� �1�R������<�@{{�L��,^�`����-\�tEf��&���I;t��~�ϟ7,�v���!�D���=w�=��F��aiaQD�MM-P=^(3�k��K�>tQw�3��RV����h����h4݊"}�eC�%��E*c�sy���-�ckn
���� J���3�&'Q�,��V��1J��Fl��Jż��|��=�t*[aW\PLv�M(��͆-�Z%tڅO}�shhm���*7ո���&I{[)��@m3����jeA��O�m����� �vn�j.C��4U����������V��Th!iA�l�}RZ��oV�:�ϗ��LA��6+��["�U3�|n�RȪ�8�X����Oalvv�GVA�ݱ]��e\����p���6��5a|~�/���rX]�3���� q�+�������	$I�3��S���F���!�F�[��)�L����K�42�L�,�� �z'�܋��(z��>#�)���8��� ��ߏ��>�U�o8��![/|�JNͯ�������C�����A�K�iW:1��+#ӈ���$ ��z'�����m��ʰrC�N�$��T7
��i��6���4�"p�9�D�ͩT"5��tyx*B�~���z�l��nA�"����0eچdQC�X�}n�)�Y�B=%:-�5�]6}�%�]+�ٰ^���Դ8LZ{��ăw��g��2łx� �����J�x���jhDoO�h.ZC>i�	��T'��4�bVqsb��\���.�)�Ю	�#-���lM˥�X�J�� =N�R6��~KC���kCW�>Ә3�Z}���z=����e�rE$�	�$R�P���^�_�����N�5׮�ĩ�W�/�P�Ԇ��E�wy� �c�n��#��K�`>�iA��t�ter1&��V\C��oj�D\��Q84��H%�K�c�A��dR����gI�g�,i�Db�\�ŧf1Z�*�&|�����6	�(cՑ�v��Rh\�մ�ꤏS,I�L���Oy�e�]�M9�,���c6Kc��$��K��g�N�h����Rƍ��X[[1�M"�l�t�&�%&��|kV�DO�&.-ӻ�~�����i%�Ű4>s�
~�+��X����nGGgv��#�pT���%l�����(#�B:����	0h�I���>�I4SP.f\�|���wp��e���yc�����>�s��.'�Լ�8a����v���k�J2�c��C���������jG2��ӧp����1����b(�J���x�u���'X�:����pk%�������YuIÕτ���_��OੇN�Z,���`jq���o��*R���rH1$�.�<g�sKe*A&��،r���EĽ� ���$d���.<�����'I�4vq�v��,��F�^YD�Պ�^Bx�
2�s�d��2g�6����X���t���8���"�����ȭm@���Z%���|^���CqA�%
������Z�P�Y�� c�� S�^�.�a���u)f�y�%���q�<2٭�5HfҒf�sA4>7��ꀛ�C�3#���>d��r�T_�����nt����ݸ4���~�oN A�9�f�,	�jeTh�O�m1g8饶�����w���������_�	�wϜ�����7��p����[Oݎ
S2�:%��F�,����)��f���*�W������=�k�/���5�vv���!��=n�0tB)��p'���h}u�C7�H���HS�D^#�����X*ii�ǯ!�<�tl�F�y�T�k0YHwQ`W��b�x��O[[S�p8*���1<��}�=�]��ٳ������"��o.����/�!�e���~����Y\�6,h������嬊�g$ҜE���
67V��hlb�P��������M.>���Ǧ�*����f��x��T��L�_]�w��l%rBI�IY�P�͛����V�P��@)�Ef3���[(E��n4�yf9de���g\���F��mٸ��v���O��B��?ʌ鶹���ì[�b �n7���n<��O��)�����o	�D�)_.JC��	��v̾���d
@�&�������Z�_���n�D����k�����B��:B���ok�iaqU���ņ�fE�#�)�sI"�A!jjg�5EA����"S�a�'<�2v�� �8甁��ő[X
�$�|�z�O���y�%��xQp�
�t6ܘZõ[��H���r��K�oI��J���b�.�!�R�Оmm�D�O.�B���V��ƍD�'16�&5��\*���G�C�-HǢ���T6���M\�>*��΁��j��c��e���㓦(�)�&6�Y\�5��5T�I�$��> �m,��j8���SH$)H-��e����у�Wu�i��:[q��$��M��y3�Q(6�.#���㢶`����W�u��{{o�`�(/1Z�!0ie�Ҫ/�� ��f4�l䰰���=����2=�y� B�/A�,IE(Oĕ���8v`@�Œ���&&�V8��Q4�Xي��w�`naIև��^������ȭg���{lJ����3�|uѭ���-�ދP���Hќ[�`xbK�a�4E�����P�(M��İ�.�CC;���m-�X ���I�L^G�Ӵl�2�
����u�A�2�e:�5��[����. �)p3���i*���\Gok O�{{w�����e�v�`R�Rk3��צ�E�*k'l�$g���]��<�w�g�,����	5���f�WD��5�&L�cٰC���5���.k�mf�C����I��-����L���ƅ�1>���� P6.�D��D��"[N�ʒ!n�f�����Y(r�Μ���<��r�t��v2٘YB�4r�au&��z^x�)��'���ES�O���?��W�Ʊ����ƾ�{�F����Uq����C4����u���E�=�H?��Ɔz=t��tw����<�^}�U�N����1�{���!'y<��ukQ��������d$횅<�26Y�M�˹���űc���`��vD�6��o�����M&$���&�R������|��9dR4��jF]� ��,�ۯ���zC�(��fSb�g�6|�+_��w��"<6fR s�Q|�{/���>R9j9-b	�����BOW'��L��[ayO4D��bU����=�T{eND˕v�o��>�;�R Y7U�4fcq��
f�\B����8����<�3���
�X����!�4�k���B{[����cH,-é��w:��5 �{���C1�5�,v��:��]�<q�z�8>���9he�ܗ��9�
J�"ss�2m��Hڝk��S����n��Kb�m&���`�<gZ�;y8��`�ƥ�e:�|'��Z�@0������}�)(݃�8����>��nLbK+#V(���I�+��Ć��R��E<�����8�������׋2��w����o~�
f�}�>��ك�S�����pcr?��{�69-"#3���^8aC��	�����N��s'q���܉����Gt��B��=�]bO�橛����HC�	���H@-��R�����Xa.�[��/M���0lGi�h��*A&D�dto���6�^�C����z7�����#��{�n���t��\�$c����pt�T^�tw�
-�7���{���%se+,)ih�{��%�N�LQ^[������2<."�n������v�i��[�s8s�:F�����J�~�^I{݊`qԡwp�4,��YUج�?�ÁU��F�.�@��l$�6�!�Da.G��rB�&VP�qR@n)on��-1N��0    IDATW}�A��9������&;�'J�
l�:�wl�{�d4pQw��86���������p�i3HZbě�.��Q��+�h �D�ǪkF���x;'���ZC��b����r#�2K��d��&%S�`zaE܆
NO� =6&aq4*�h҅TYd�~��@e����:�Vd�)�&gW$L.���`F1W�z��C܉��UiB	[G2�F��#��1����|�[Y��S�!�q�-�֌�fNY�� "df",i '@ؿE8L%�ؿ�C;:�%��t�,S���Z����֢L6�yW��hP�IC�o�Z..�$�����#���vw

H��eG��1��t-s�b�#�c���Els�:��gg/|~�ei���%\�>�~C�4�:;<��v?�E_YY���PkS�(�L/���W��J8��^�8�d�6��@�հ�"ݦ�яޮFt�7H��3�V�;`*���ʗ�x!�	�q��4,.G�ڒ͠�0،Z�����P%�.�O��&���L�J��E���pt�_�b��ٞb�p�h���p׮ݒ�Ng�}h�w��Ή��O��y�-X��Fz��\3�����2|v���A�
�ςH����G1<>�X� ����`D!L�}��
�t/�������e+��f���r#��,�Rv��̈ ��#)Ye8�N	��f�7����@�|�.����a	�S^��~y~!*VV
HF6��шG�>�����5x\4�6��j$�S��qyde�G(���Z'&�	��5r��TC��ɤ��,�Y,��QJ�Q�p�[�>��5q9��b��gm:p;0���4�:�kj�5��Ť�xG�-�@.5��hM��x�O���+i҈J<dCd�F�@�o�SDP*���I�cgN����l��1(��/ـs����*�__:F�Wŧ��0>����-$tԼ������ݿ���:��[p��c8q�=օ��5?����	��o���{6eZ1/�<Q�,mGu�A��5����8��Ȇd�>}Z>�[����ԟx]n���`"� A/�ך�_kv�<Gy
���4_�C8�/|����c�����?��_�*����S���!t���㢓�q���jj�A{�^ܘY�_��
�>se�UE��E6����~y�\��(�!�K݋�|�[�C�~��fQCKk>�O���E]�# P,�%��5Nɾ`p�@SC��}�-�������ׇ��f4Ndl-�c��i����r�`g:�hDjY����F��^��5���i"����!�Arn
��J��;�⎤�E��+��t�����e4�@���Z��O�b!�����6�	��sH��b���̭����TF�CE¯�R�U
ԏUPd�E����)^,�9q�yfsB`Z�����7�h^�!8v�F�cZ����E���e���Z&��d����#���4�_-�ȧ����{}��������_�EmG����������V����:���V�3�;{B��e:���I���Y\��Ս���Z�^�S1Q�?���8��^��֦f<x���4B^��<*D$-e9�,pN]���^����C����!��,"xB�:�E����&n����3o#�2	�� ��Q9�y �8��^����D[k3C!�4գ��G��¡C{DD4�0�x���w2?�!cL�0;v�X���đ�a/���,�
q��
n��D�!G��}�XtS��G:�siI�o�u����䩱Xf(��k����XZKb+Aj��f��$5i�����ӏH2+�+'"���S\�.d��t�b[K����@ۚ�j.H�EI"�5�TtUn".@��6�_:s��ǆ@�w�bL��܊��;`��s:�&�������yq�r4����觞��eǍ[�Pl*�����L���&f]☎(�!��M�p�\��V2��
�۹�5��f�����jb�Q�Ru�4׹$��|d�u3۰��p��hW�`����S�ÊT:+HBc��\
�t��-�nA�[Dk@>����������El�X4�r������ػ�]M����P͈gRиx[�X��06����5D"9��Ɔ,���i�*c�+%g����I-iy$�����ݞ4>���Q��Lg�<�b#�|6�E���`o3�W�+1�[���Fn��x�ǡ��YB��(LW�aX��@Ew7N[4�GF1?;���:��&��|�,�R��\�D&kԨ��k��Gv��QA!�����"���16�Y�'����Ī���&T"������*��	�at-�^�w��% 7�J��ur�s�M�3UԐ,�qk~c3��������<�E�={f��0�  ��"V5��$۲��qY��ز�z����NVrn~�fݛ����%��*�q/�U˲$��؉F�����^�z�o�������\K�9 f�������>�XNy�<]��UU�+G�j��ƺ���b�#h^qw�@6�hx����H��qu��Á�h[�4�ֱ��%`_:��8-�j���e�N?~N��8 �mau�'�0?� ��oQ25Y|&V�vqebs�Q��0՗֟��ZU�+f����R\.�1�ׁ�'G򐎙�K�VO&se9�9Xn���g�8=h:��-e��6��XO��^�4
���7,��Z&֊��\�<_�p�9:$.�Ԅy��r;6w�x��C`xZ���Pf^��|R*e
�Z���ޱ��t�{�I�!�1���NU��D��㿛�V$�����H����̈́�\������>|O,����X�s�M�$݇�r�z����ɜd�7�=���i,x�����=�GkSH�^:/r�ܟ
H&b@&I���
�X�F�:�*��]V���߉����a�'�2�"O<�,��/�;�V�܃���f�߇t*#V��s�H$�b@�����H#����b�X�e�x�o}��N��]f�����5��:�笀w�~誱4��n��6ߜ��۠��kED�Ik��y�	�����'1�/�F���Ǟ��¼�b<t�����9V��ft����q;�b_�)]sk;��}����o��x���(jttt"�ˈȷ�����r=�!`eP& 	���͇���p�Y)������g����7��,��׹��Tzz���<�T��(�wd7�W�i���_8�/}�2-�t��I�[+c/�r��y�ݰ�c�T-�VHWT@ �x�֫��P ����%�3i���#%��'���ȴ@��<Z�����҂�o�Fs36���۬�x`���KX����~�2l;I4���)�5T��)}��Z���J��Q�� ��M�M��9��M�>��M�~6&��6��>Ԛ��KG����w��^�xu������o`i'��WU�'V�E�A+U�(UU�1s��rz����O������0���׆��ϼ�����W���l�ۻ{�z��;p��w�#D��nn����Kx�Wg1����߰����䱛𶷽�'Fq��y47�q��M800(�˰� ��@�h��(~}q�,�e�O��%�5�Pr�u�6�X��.���^?��їPOn :��8v���yn��W�����EKs^��{�9�{�x
��~�|^x�y�}�<��a��1&����N��7�`(,�>��iJzo��3ʕ���L�䡠ƕ.q?X[ݐ��)���0*
�2I%�<v�P��.Ҷtjq��N`ayۉ<.�΢\�-�.�q,�9��7w�f�"ǿ��ȗ,� �Ak{n;Q��\6��97���*t-��44�O_���a�S<U�tLaS�1���]B40��`B���G8�	���$�Q�`�\�� ����pelR��8!�����H��MhD�\4F�\"fa+.!^mE5���W��(�#{S�g��9~f��m��^�����%�� �ӹq�l���?�d����FM#M��i�t�Z��_�u��Ў�{��!�m���)�&��x����u\_�v�&���&��D�8q` {��ඔ��6��b�C�⒆���2��-"������T�FV�&Xhv�����W�Y	M�i�����#��S��RPJz�1��zc�<{[�
�VE� G��Z��r:m �[䫯�������)$�8{{:1��=a�4�%4�AA���V���$"x8��:t��`���'c<S��j
�M
m�����$���-� *����Tkr���(�.#]Ա������X�J�fw�����")5� ��W�#�nG�BuN��7�Ǳ�0��L�� \�nE�X��m��_���k��G�=-s%�]<q�׬
/��Lɸ&Y��9e�Ih��ƽ㍷K�5QX�W��<�6iܘ[��VT����[$P/rK·�^����?�p��Y�[��-HS������hmk��D�-#͆���M΋n�y�]���p����:�~�t1�o���#8u|^��
�n�:jQ8� E�\���K�:��+�t�<�>���|�׸t}.�`��i��^R���X��JI�9y���KgPQJh$</�^3��L�^�:�WF�ETnp�@Ђ�1fO��IZV��W�be7�}�@a�7����녟��c�7�&��Z A�Y�H�(A����:>�B��4�����yfހ����JM��*���; ֤�ڴ'5ir�~I݀N1=��r	m-M"J�t��C�"�hwg�T6�Ns�M���@��\�2r�8�Z~�=���ɤ�9t�z�ٳ���"��MH���a��ǝg�H�)2�����҈e�9��c��4��>MN��`#��z-҅8��� ��T:��F�������(�L��I��2Ch6��� �a��4����'���&���3X]]�07��ׇ����N47�i�s!��}EZZ��aj~�����/���A��B1���Z�\x����g>��9�i�_�8��}�a���m����6���Ͼ��p�� ��.�CX�����U#@j.�t�v�_�!�f���bŹsW���_/�-���GO��SC�ni���F�ˎ`�WU��5��!�H�]-�cN��L�RA깞�Nx,:vQI%j��Yg-��{@@��X�ޫב&5��D�5��U�n<��J	��~��;e���mѱ;1��W�T!����\Ar�X�����cс��K� l�����Ks�
�
�S�n�TI�(��Z�(���w�ZN�;��%����0:/����!����4F�sW�V+�^L��>v�S���g~�����_��n�z&��&x_o'�Go[��vb�?BGU�y��-������!��`ycs�KȤ�hk�`��N�U�ae�w�5�'r00����_Y��lK%�u�$Y��:ڰz�al��2�t{�J�ޜ����ؘ��
�̉���אLa�Bn�>�Ve�����Ǜ�p
���x������ ��,ҶH�Ѕ2�"Ξ=/�E[����f���%�)v�E
�L�W�P��������s��cJ��6�V�nɦv���̗��+Xߊcbjk��6�X\��X�7{��Q8}-���ԎtcD_՜r���`s@�9�ÂB.�f�b�S�!(m��RM����������,@�fQ��B
㎩�hxY��!;�3��Цi�*t�`�>o�ע�&�&��}�Ň?� ��\�T\k���
�t1i4n���S�2֧�s^������n�&�'�LÆ�_�f@�p~g�E)Ď�Ş�&�]6T�(J�����v�=K�Hdi9HW{#D�"�ݰ��J�C���=�"���c��Q���|��x���6��p���ZEgK@������"5.�΂�RR�ay7���\�X��r��##]6��G�܀(8��W-����Fe_��=����ge���65��6P��2���^�Z����߃PRan�ž�6�_�(T*�n�191��5fl�u�-5D���#�fP�����ʼ�l�JȦw䙥�fu����(SK;�]�n*�L6�VDww�vC{[�Ҍꁝ��h+(5d�6l%˸:��˓�!����DGCTT��< lB%`3V+gE��е[�����
P�^I�E[?�H��kӸ��2qK�8��Y�&Q��E�t��@�q�X8x�7�X�ZM�Q���{1���a�Ņ��a+����9�^����p��4���xl�@���,J�2
�2��e����U�./"�A_/*�t:zխ�Y������9�l��,���#���S(zB��4n?1�7�>�N�ȜX�9],Bh�W�Zt�_�Jck;.c,�(f޿��Mp���B,V�K/_���)9Dm.����dY,viR'Q�Ġ׳��Λq|'�6.�h�`��2M8]JdK�\�F�F�<�2��]EDܻ�c�-��0��s�7p��4�m��k�J��c��g��e�G&�X%��ј�(����R��Q�6�?��攀A�����fC���ϯ���*NR���Ig�zM&��.._|�(l�M��9��'wQϧ���c��&�4�ɡ�W�NK�����>����6��ٓ�<���C���jj˴}_���/66�8[\Y��2�'�Ż��eym�aQ>���,���@� D-���˹�Hv�>).��~�d#��n�B���r�.����p� [5e+��E�@V#��Z+�P3@�(����6�pz������G��Iݹ|e_������kp���;���6���c����;��e�����}�a���!S(�v��N!�Ӊ�|�x��߉ps@���nLBN;Z��ȉ�E�ynGҀQS���kF�Zr��_�������ʵ1)ֹ�v:u������"Z	m�>;�ݵ&M4A�2A�_�Zxݻ:��'���bb�lv�I"u��!�m�&�A�"Y�J��Mg$՘���+{���@+�躵�%��ő���d�P���n�{>)���	Ҁt��/U�՚h^�^7JBu�>�7k������==�>
��c�[x��I����^���9P�(s��U���4��t�����ۏ�|�����VM��˳�������;i�E�6*��D^������#�+����Z̃�g�]�%ːd̩���tE��y� �e]��^�Z1��Ǔ�Oa|>���u�'Gk�=�+�="X4��UE9����/ �4�J�:3�6D�>r&��9h#"��M������ܧph����B����Ol>�$�)�"f����	���
8x�0N�|���L���RǾ}{���ӆ�v6qG {Î�ְ��+�F���*c��n�v��T�˫؎��-h����#�I�Ӎ�e�M���mA��Q�Z���HN���� �"/����Vo�*��-����l�Ϡ�D-�˨�a�P�o����VL�Z�H%��Q7Nk������M�o�
5B��C���P��anmDQ�����ӆ�ۏ��<A?F''��(v"��vc��c:��Eu�ǚ�!v��Ў�R�]��81(��OC��ڑ��$P�,��2�N.{��qpoZ��bZ��͎f ��bfq���	�����zV���R�Bv��ְ�m��@��6fD�X��p"_�19��_��RL|޹.9��l����nF��
'��Hȕ��nՂ�Tӫ��\��fV�)�h���{!�1����%���K���0�ۆc�a��^�[�����q��B��kbٹ�(�J]��e�59q�@?��D���i�g.���
&'�����B���'oFWG�L*�Ud���I�R��r1#�,�RjV�EsLd�_A<��(�R>)S��G�q��C��O�8�qʔK3�SG�jC�����y��:�D��/��P�sD�')6ጲ3��7��V?^w��K��Qc��i��V��ynEi��6�2�KT+',�6�i��y�a!�_< ��CV�d9�:������6�rdH&�*��X�H7���.2�w���p�ll�cn~Z��{���R(K�7m�3�2�����]���    IDATmB�����jŵK��^�n�"'�dUЫ�T��������x�-�s�W��I*G�U��el(���F'f���I��ʲ4o>y#���#������O#�,�v�WJ�-�%d�b�{�mG0��Ex���!�4`�|U v�9i��X��@wx�!�R&6�04�9�x��,�̉ ��Y��4���"� 4����{LD��͇i|�ߥ �TD���l~��Zy.�iKCXlNȁ�{
��r�8���6:�5���t��� �!������w�%��ڕK؍��n��dCP�e$k�Ω�P�y�Y��dP��nG|�=x��C__��N�~������T5�N�K�9Jf(d^�@�d���(Ia��d��GiH��/
h�Lq_u��*��HA=�X��<��DZL��2M��/H4MG��K��[���nX6�>p���SY1p�=�&Pc��ּ��y�Z�V��A5�x]2��{�x��@8Ԅ`�I�ǳs�x���cqm/Cr�;kh���~�x����)H�ʸ6:���oቧ����9B��G�X�[�}#��>���}����s�_���hdd��v"���19���zF�Xk(���x��w���W�L�?zO��E��9�S�W
Ջ�	�HW;��<\�-t��pW4X8)���������mB#�=cC���a���5$�W�<��(�`�v���D��"ת�B��@��$R��8goX��nC��S4�BQ 2�����xLjjd�4��)}�M����󒅿2`�V��=�!�Z�rU�E�p"�����#�Qh��X4�_����Ϗc7��bs!G�:m`I�yܘ��aC`���[����'����>�[�|�g{��_��ŝě���1-��j��ӊV�{�;1�ߏ�������D�Y.s�J�����F,���U�2t��#��΋�f�9ѝ�l���m���K�ߨ�ji��b��X�6�=����S�AGu�Cv�-EL��cP�]U��j:�f� �FÎpk�z:%�7�ؖ���������x�G������.=z�p�qp3&���h�$ǘylE㘙��B��⾁A�t�MH�bX^^D.��ͷ�"�0�6���)�#n��r�����>�N%�m���;N��j'����<����܁��v,,mblb�3�_ڀ��g��v�cm'%�x�P�D�+ڐe�IcP��-�V(ccf	s�^�P+%�٭�V�P�������g�*�Re���@>h�`����f�n'|�7MV$b	�<�� |��I���%�|n~^�Da�$=E!5��!�/sJ �3��PS|'E~�!0G����ޫ�-�D�j�uX�����n�i�5g���Eй�8k6�6��0��2q�R8�~��i��	�q��=�
�TnC�*�Nl�c3�x��E̬���ElJ�GgX
�}]ax�
L�6��dU�v�&	�W�汽C6�::4)[X
��Z�y�rC�I�T�RB��@O{��:��'���*A~l(�����0��0>'(y��hW�?:�+M�ӡڒ����&�S+�f�ߡS�D�a?���>4S�M�1��s���%�K��� 8C��F�7qe|NRk��Jꖒ���w�@[�)�������"L'А�/^���K�H�i��i&�tҫ��]��D��K�]�e=}�n9���Y0��,�kH�ʈ�s�_��ձ9l%
��-�D�`1LA<�2�@j�6�vHq��N'HWr�j��7��+���~7�>˰5�\��t��i7,�l���Ʌ,�.`jjRF�tu�n��&c<Q��iL-���psHh l��&titS��H�	򨃔��
�#�R�+��8�L
��8s��V��V���D(j�%�~3��׍�I�& ¦�����f�JE�fG2�����oLc'��4ךn:7�PS��കpx�G	���E��ҍ"K��o�R�<��k(Y�2!`�#����fI�nXx�{��	(�d�+�D�)�l
�יȼY��y�ŭ���ee{)Emc�mR�^�G�W���J
�FSi�G"��}Jօr12~?�5�m���yM�Ś�Թ:V+��(&�ǑL���Ag��G��J	:��Ւ8��:rP���$����|胿'�w�E�~�������%�(������/)���C�7�?�"�������sE�������NTR8iɼ�{l4mfC��3x��7�4���hU5aJ�&5�! ���/�j��72$�.��lP7����4�dC`��0;�[�^4Vl�4�Y*�D��\l��P,a#�Z�'��J����:�N|�#�?��b�AЈ�s�/�_��M<���p{<8q�A�nL�����/��7���O>��<��Ʈ�{=}�|�ӟ�������=�0&&&�ͧq���O>�_12t?�����o}�+Qq,$[í��.g��u�PG3ڬ54�3�p�`��0j�>/j��>&O����� ��+{ufc��0�tF#��֞@��l^%���݆���	U�6�s�r���,�l
;�Ԟ�$��1�4y]<��Ə{iT�z�	LЉR��4(i��eC A�bP���	��9*҆��}p�|��g����iL�&Pѽ��t�I���B`QQ�U�!R	��f�˷9�ɧ�����V5߽8��7��^�Z����M�NQ|sL�Hs�MG��B�ߋ��vq���+h�"�1ar�BMH�rXZ\�n���%�/� ju8\����1�p��
���������J�J<D��A$Sv�%N��#��߁�k���sO"�I���Y&
�u#%Gv�z�H�؝Q���@��n��>�[������]Sc�H�X�Q�J.�����/בL01>���5����;�o�>X���]	=��SBb����8��k7�H���ݐ<v��뫢O��w�[����M\�2���8��6q#�-�26���Mܘ^��N�@�����#�"Z-Rl�Ɏ�b�'�n��E8ɼ�b[s+X���VL��
�J�Fd� �F_�������a7��(��-����qRzȏ+����ڼZ��ΣN?d��.<s3������sc}s�ݴ|fA��;���e����@&Dj�U�]Ù��`4���@ ��?���l�4��)�:z�B88ЉވG8��V���o~�����݄��]å��YN��9qC!ǰX�o��Տ��fi�`�\v���Ai�$�{bn	Ϟ����� �llZ=mM8q`/��#8��X��`7`w���7��Wbx��$����E$�S-��Dv��4�,�*�,\�a?:���4)u�a�\��B���LO>	��k�\A�9Q\X)f�	�i��G�D���E,���n�qDc����'�B6KU��#��I3�Z�`��z�)�y)H�����M���Y)�-���W���h�]�8�mMAi�
��4#�jv�e=��5)L�t�;�G+�k��,��ͥP�{F.�^�mG�q����2}�����wMe��0�M�ܥq̮D��]p�!�S��8�<`���
�)N�x4��J�-�A\KF�����ێ�'Bs�#dD��?lt�kN}�%��m�I����L9[[�p��wc��KZ�<6��\�ݘxm��H��L�$=��+�XX��T#�����#6��t({�*Ŭ`����߆;����ఫ��\�#��#G�G����.\��	��NG�JG���t��	�Ҫ�P*�$tmfaۻ	.Z�e��烳�"*��:�i���0�6�$Es�l�X�/�O������V��؜�Ś]��p?`�b
~y̂�L�IGT���W]}���Wѿ�1�=Lj��b-S�BAM��2��kMj�9}�F�P9.B됴aUD�X"��i����1݅hy+�g#dޤxr͙{�4f�y�ei�Ѫ2���k��g���� �J���a%͌C!�+�<�lj���>�>����@gGg�=�������[1Y�<��PN>>;}�ϣ�&��7T���+Ey^)�e$׎�皲�pTM��L��F�rT����❮��ޱ ��V`��V�uI�j�t%gAǦ�ֹ���Uc��,��Q�J3FGU5���4M� �J�n(m'5�._Pi�i$��t�� ����Z��!x��g���~���%؝��u����=���B�^�?�~7�x�	|��_��R6���8���˿���0���/�����>��f��a�������W����!�@�\�>�������A/���x�&KF��n�F<4Q)fs{C�#�%b�e��ڂ��X�y�ז�\Z��iC�Z*�W������8�1�N�k0��j~�9#�BlЙ?�hЄ�W�#��	��M��H?���FѡE#kA�k��P6�V��ۅA�`��vt9	��l�]8;����M���b����ZP5�H �a/6�I���Ttu�ԑ�O=����5!��׍�<��{��د�>QӃVo EڼQtS+��[��ڊ�f	{��\�n|YP�hq뱛p�-7c'����G$����U��T�!�Q������V��</���#)�ұ�p%r�w,v8����~�]H,��쓿@tu
��3������H�z�w8��=ݰhl�lH��_~�s��ԭ��r�����˯�sA{W�x$�+�M��œ(x`�1uc7��UB�Mm�p���ر#�7��h?�0�]�.�5~"<��w�d����%"T�>t�{���L�����bl|�NOW旷���������2�ַ��=�=C�`�6��%Qk�2�<*L���8��^��@>G{C+�R;�kX��@-�K-�Z��S6��V�?9t�tZ��h�͑�]��-Ɔ��/O���Qm��y�#U����ێ�]�/</V7��y���;r���߀����Mᗊ����k�����(�Y�u&���Ex��(�5�]-������˶�,n<@se�܆�J���Wqybe�2KC�R�i�ǀ+�K�"�Y���$ٗ�,��I�U]Ǎ�U<aK�EI2�Zj�t�'���.�8Q�V�m�!�[VdJ���.^|�F'�asx_}�X��Ƃh��l1���ي�H3�ۚ�) բţ}��]�(]��?��EL-m#[�A��h��Z�¨gpdd��c�NY��\	kIܘY�v� �w�����8�pw˱�h	Zu�R� �//��&9դ�!�߈��+Ӹ4:+�Dr�lZ-!�8<��� �+|C�?Qu���"_�Å���dP'M7�!P4D�v+�$*EحUXk�me�rx?�8q�$������(kp|H��Ϗ���[�Ҭ�u�4�����P�aO)6���D�
��C�3��<5dQxlU?�_,p{ښ��(��ҝ�"I��ʘ��D`'�Ƶ�Q�|�Z�M�ݷ�C=]�K����ړ��l�yֹ�5L/l��$�J)@s���6�4�i��Ui>Ģ�T}C�e�ءh�<F�()',v���uDw��J������D^r�=>�ʖ��&a8Ծ�zĊ�����&v�)褫؝�w,����@%������!�dաiE�ҹ]v����rO�0�����L�H�`C�� �],֤�&�����M����4��NL����7�@5f�b
��I��T!�n�8�-�)L�[��I��\/.��:��Q��?e��o6��)2���5�����J�\�:�)+��鰢%B"��/����*<�І�h�!p2��-�4<�lT�%d�1��|������ކ��&�eaj�Kc���:&nL��16|$L+TS�mo�a28�e�����sr��{�}=��XR�I�cW�B�ٸol:vJ���5�����(?_5�j��h3MZcU�Kڤq&p�,�U5�}Z�Sc��!y�rOc�B@����dA���i�j�"V N�u	�$�A�>Ț����=����|��#0�-�g?����q�긤;H=A�5�������×��O�@/q��-����7���E|�k_S��l�����_`p`��?���}J�r���xum;w�#b�����Mm^�Ji��:$�F�\��t!w@&I�lJ�H�Zh�Nǝ\۫˨��� e���Uq253j�d��55�3^W��4q����=�F�RQ�:�9E����'j>%"��Qڨj�#\�8��	��n�Qa�
�����Ձ��~4��3�禗��i\Z^�B,�T����t��dt�f��iiOt4�ѥ��������G>�����/~�&|3_~f��_�֏��O�XCM�3���A*�����w�������W��6#�N~����r3�����򕋈nn��[O����*���ؗ>亠�u�钆��7���?�ո���|rh�����
ɃV�f)�)�����a���83�2�Ņ]X,E�ZI�Y�-S@jw�E�_*�%��}��.����uZeBp��E�n�<�p� �L��M��N�a6��p��(���`�4`��}����ؿP�l�/\�#�<"	%	����E:>>*���Ȱxs��74�w��]��f���1Vע��?�x�$��wX����Ģ�k�����ٱ��D��<u
���%��8%��l�jY�U$W6�6;�Rb(1��Թ�2�Pč�,&8�'�BgA��$�T!�\�,�fW^*�j� �)^cC�s�L<?旗��s3f3P%�&>�
��P/5��tܐ1��H��kx�e6�$l�O�k�y� 2�4�.�4tЉ��l��A��F�I�Pډ��:�勸1�&����E���p�t��b3tb_;F:�b#�i�$Hk��@��.m���l�V�!pU�\]���ώ��q�� �j�����t�1�ڎ��]���u�άBMg
�� �#�LU(����>t���n;��Y8݁B݊�DO�xI��d��C�dI�W3�i���'�N�H�I�K�6:���eѲ�Wh-:�����h�p����*5䎲�v�b����95/�ps�1<q3+QT,N9���M$�5��f�+�������y�,5�\�Ն�63+1L/mbq#�T���8�P<h1l��hrW�p��pZ��u�e���!�I~l��3��½�llϽt�O�uc���л�eb1��4�\�C6<��lT����Z�	�����]jz�B[�R"�R�F���E"�UD�el��������
���{��ގV�%gZ6iXe��*�G�t��\vqr�46+�m;tsх���*
���Ng����b�#�w��[nB_O@lS���=��R|�������z��)�l'�M��F�[�t��~���as�aw��f<��c�#]:*�3g�K��<�����80B5���b�g�*�\�#S�!��blnc3+�g�B�����#�HD,�/�8U�o�G���'� �����8�~������3E�f�n"Ȧ�P@��������6iD�qHM�UEI���B̀9Qc���L�M�	b��b�T��6�U��Ё��� ���t��J
�K/����:|?v��J��d��HgT*-�&��?�BS����~�=����]�^�4]�.]���
����Y����J��'��oUy�,5v�gΉ�餣��b���'I��(��s*�#��aeuKkt+ʡ�hE��t��� R�x�%�J\�j"��������)�kf��CuNYZӪ�SE��_�T�r	o@����&D9Ԫ����!���)6�k��i�������AW4 ����'�����.^E2��Ɠ�5Ҍ��y|����P�+_���|�n�;�/���q��!|�K_¿��6��)=y_�c��������1q��vڢ�V����ƙ#�WQ�X��N?��<R{i�L��Ep�,	�Lx��'i7���\n�=�0ܚ���ui6뜢p��^(�j��fJ:�F�����������I���׉�T�?� ��/�Pu@C��1�f��4l,�1(�B��Z g�z8���^Dat�a���G/\�������W��U�vN88��c���f�8iܕ,J���]'�|�ѿX㕆    IDAT���V5uǏ.�����g���)y��m(Y-�ۈ�%%?�^��Z~Álz�X����D���Gុ����+K˸�����$؇��<����T=�����[���~��Vw7O�x�s,Hq7�����GE	n��hqZ�4uӣ��:�vam��bo(�B��U8�DZ���Q.fqhd���qӁ!��yLN�!���L!�������'G-�.*��T������t� �����b5������g?}��կ$ ����-S 8@ǿ׮]���S����U��]xǻ~�]}x���pcf�`�ݏ����܋�����,�5�����'ʝtZB�(��9}e�x�*Z�l�0�kHml#�4���&jE�!`~CVh4�M��(�Ħa��͍O��PNJ%*�)?�+�Ft��+b���@���p���7������Ej��T\��h[�����%�!m�p��8��A�L�@н���~�^�5�ֈ�0B���#���_�?�V%�f�5���צ�x��_cv9
�p#��b�紆��r~�a{��oOA/زh(�bC�.U���Չ%̬f��KV��k���f�PVn=2�=s���P�L=�l�2BY�6��b�e�&�����æ�,�����=G���fw���h���R^l
Oi��ӓ���Zނf�
M�W���R�p�� <vH�͵H����^x�*��9��؈�j�bVɧ%���3�HS�pP>�V!u�ߋ�5qz`*3u��-`#����.*5�O{�ˀ�Z�,���49`��E�+;�`7[���2�O3�/SНFg���8)U��9�%qb:����~t���Պ(�7Ft�M/{&�����KX�eP�8��F���4t�j䨨S�dD<װ��T2f�ci��,e�u�����)���C&.���τz�X��*�$�Y����YL�O������N쉰P��Vd�f�EA�j`�̮��\�����
�w�H�JpR���O틙�M
F��fPͧ�����'�o�v�(�\��ܦ�+�f���UL/mIA*�Q9�Ȥ�cA2ʞ�JڌM��L.&��JwC�5h0QD)CG��y�=�0e��t|K�dyH}~Tk���u\����9q�bv�R�!�} (�2a;'��q2�v�3b�K���ߤ���5����|=���t�p7��r^i�̟e����6��q���#?\4h�� �,�ޤ�Q%Vf����)n;kWixh�)�V�ü:�1���cm���f��1�*��	�>����8�Z.�b:-|mK�*�!B���8��wߋ�ϛ�o_JE�qJ�US�*��L�kO��<Hh��P����W���'�'?'��j��Ns��3��rQ���R�MyՂ��(�~�9<��_c;���*wFN��h��k�Y1r�*��f� �#�$�: �e��J&�#J��ƃ,
[�3W-׃I��A}������&|���9a"�q�P�J�BA7�t�����!�P>4�8w�e|�1��"{O�Z���ui�~�wކO|�c21x衇��g#�����7���$G��������~]�7>[��~>�'��޽���W��Ǐ�~�&]�`�
�{:�޷�	LBڝ��+EĮ#d�Ò/�V$�a�M-�]�A�OѾ�%��1	$����B�x\�Qg�"\�oj�_�+�g��V�Z��2<L�v���2Ǆ� �	���Ȓ�� C�Y*l�${��↽*ݷd��u�;��R�ӭ��Bٰ"л��6��"�ׇ���_��O_���|i݁Dł����BɪK�	�#�MNK̆@�VQ%�]L��s��O��/>��oUC��K[��������܇�@+���퉬)g��t��%5��9�� �#���؁�����𝇿���9���o�]����i;��_cq0Ά�ŁsW�񝟞�����U��Ƀ'\ݐ	A]����O�^��V?v7�1;qk�㨥��������ZXD߬��m
�r؅����+���p Kk�x��XY]���D�[��˘��~�+X]��Pd�x�,=�Q�����D	�s��fp��9�'�h��>��X�@?y򸈏�6@~���n��4�tϽ�[X�<����t#����؊����>�مuqL9|�F�Sy$���p�K�kkHAme��K:��n��2�m��΢��!�T�q:���h�T����D*�8���R�����(7c�%}I�>>Pr��a![`�f}�o�{?��2�0'q����ϗ��/6f�Xc�ȵ h?��|�t^c��?��!S�g����p���O�HW�#䴢�Ń�Mhy% �16,.b�*�7�=?���<�͝(�X�1�Ԟ��I�����v<�Z^R �q�.D�z;�ù�70�D1��LJ9%|N]�GO�<�����">�tk`�U(հ��J͕�u$�5�K�,'G�.8BZ�QTO=��^]�.�vrma�P�X��ᔰ���D���3˘Y�#]Ԡ^u��ޗ3�Z����0��袡Id<��[;i\�6����%#C��_'hK�RNp�݂H��}=�ӥ2*YA���ށxU�R4�W�永�@"S�]��5����ky��r*y:;Zdr �Rp�*�Uo���x� ���p�°'��Ws�9���ΰ�N@W$((!7tRlt��L	�N�0|7W���s`�B�L���|v� k�X��:-�Pʧa��?���C�D��1���~�P�2ټh���QḼ`|f
��$::[q��C��B�n�VIK"��j�ՠ���f��__��/\DZ��~T�6�Dq�� B�ڐ��H��\^CC�Ê�8<�%�"m:s�����ƕ9��i�ZG��u_��l��U���h�7]�8��	��r"�L��as�a� [GG�o}�)�4b~�A�`B!/�gn�v��dY4$g/�a7WS9jq�<p��϶)��,�Mߜ*�}l� AĽ�@�����#�M�l"���6��@MT�*�Hi*����������	 �҂$� +�
�y�8S�����uռ�!P?�a����!�2d�'x+�ɮ���ͦ<㤔�x�Υ�.J�������?�t$��ӥ���߉�}�hk�K�@�=9�<ӕY�o>Ol�mB�20'W�PJd��x��S {�*ֈ6��HR��Z��D��^	�g�
�;����=�09Y ]��y,"y���_�lB î�f���w�w��V�v�&��T�g�M�q2��ƫqޑ���
��MGcm����4����Ib6S�%^� CNI������!4(^�n [.���x��"��I A�K�.�X(�ԩSx�����!��O~(@���Ɖ�O���CϞ^|��ÿ����w�)�p�uw�����>���9|�arz�\A�Hs��to���mV��L��4�Ztz&�Ӗ|Nr�+e�6���j��ކ��[ص:�6.�u(�3rVqz@	s.x�����RVV��	����f5%��$�f�ƎBB��Ui��tZA�5A&�R6�fSF�U�7j��T���%���	ks3����<4��˃+K[�����E����V_3
�U�u�K��=T�觨�e�q��v��s��G����?�[�|�����o}mv#q�'�{ $�,�t�kL��x:=�keAuY@��u��-G�7�?��c}mw��N�r���!:��NrS5i�_�Q��Vg�:�u��Xl���'c� �7\�vK�
�����q�\��bb�Զ$��,8�mxN��Hʩ8�~�gn;����N<4�xb3���*^������"l}m�|^OH��D*�d:���i:8�e3�hPPu�����+X_ߔ��)5##C8xhmA����Ii<����#�܆��y/_Gk�^���nkN|��O�W/\@Mw�gϠ4	8ϕ�+�Q���ؐU�8mJ��p;�}ri�U�$�7�>;�r**(�P��3k�lŝYPz6
�'/��pM�ł����#��(�R6p�,4�Ҵ�q���ɂ�3��w?p��WV��j��@��!��b�!��k��X�MC�j�������B��W��Xԑ/f�s[%Dlog3��=�tx�M@�����`']�j4���Mcqm��XA��ڑy�r����12؅&�Ulp��+�t�܌e��+c�^J���R	���X�ED�n������<<H�R|s�N�~rg��Y\^\��N�,���ȁ5�ቨ[��D��;�t�����C{��2�|j�y��Hayc�Ӌ�Y�F�b���*"D����8yx?�"!xi&������D���$m��*�u8�)���˹Z��a��`x��Mn�(��%����6vp}v�+Q��5XXR�I�F�"J)��铤^�׀æheb\�)AM��z�L`bz��怲Ŭq_S��]g\`��X�lǑ�>�%��Yy��=�h�0�:6���%��^���CRl�aP��Z��&E%��U�x��$3�ɮ����G�(�ZHȄ��B�n�L�R���Ņ��<^�>���9q���4�v����8��.+��,z6�Sh	5z��NIs~���y�22e�l���<Z�卜:Q|,.PE&ǔ��e�4���(.�:�sb7\�Cr2�K!�Ս�ՐÙf���M����<�ץ���}px��Mdd߭�֐��|W}�!��t����F��LZ��,��N��.���kS���B���?	�X�ˁ|A�)T��M34)C�w���?��Q�Wh�IR�&��`����q tN=���*�	T��B�mR�(�������-g�#N@�
�bE}i��`b62;%�B��w;���4b��vv�uy��g������t�).�4J�4G04\���I�/�U��-�����{���،��@]���8%�I�;�il
��C�Ah"|6%����2t�ө��Ԑ)���*�A������B�������#��M�����|��QW?KC(�(�8vt��ԃ���M��)�$�*i^Ho�{4�i��F���{5�2�Vnz԰�ɛo�#�'�'k�H�f�Jn]�(�t
K+�H%3X67������2R��ؚ��/뉍��䤸%B{W�����5\}��ͧ��ۍ�G��#Ҏh4�������fg�J�1��z���M���mkkׯ#:=�*S���3Z���nB�	�-�X`��+��А���"vE���J�PR#)�e%����<!��gE96��ƓBa	��������7Y$܏9!P?Z�$%Y�����I��S���Uؐqbn�wO�FB�`lu�����-"g� ���	�d� ]��hs��� �h�x�{+!��45�}�:�sw�z����O�V5��ԯ���?�[۹ʭVw�K%�L����:��e졂�*r�݆!�z1�3��ě�p^|�E�<p {��"�P�rN�$؜t�HƎWƢx��g1���v8|-���K�&`"��T�.����||��W�]��q8�T���0S�x:#�͆�Ca���7�o}�.��.n�N���+p{t��KwLG!���N/�B-�y��pƒ)\�zW�^��N��`�'����șT� ����G$��������������҉�=�_���r�@=���-|��?��nvw�{�o�F���I�2�jN����M�U]���J*���l�Ϣ�	a*6����*gI {
��P�X�s�B�"J0�࡭d;R���Do�.�?}oyϻD���C�.�!�07~D�v�ߏ�� ��Ϧ6]���!��	���!�D��'���j�=�
iq��׉{;�t�C>�]m6,`8!���2!�2���h��.T*TA�1FE�������� �7���Q��dS�X�"H^���s/^��|n_+<D��y�V��8��u�8�{{#"�#�;�)��2&6v���I,�F�����KN݁V)	��7ľ��Z=�j����g��C��y�$V7��ϖQ�y��"�FJ �S���8rp��1���#��cay�&f��̣��D�*����Rϒ�%�Imi��	M~�n�"�3�;hyL���\ܐ@>�;�1iv�P��4:���i.����r�ŔnКӅ�TW��qy|ۻXlXlnE�euK�b
�\�=-��u'��ύ�vFP{N�2���]����]���4N6gP���b�����k��2�J��[��BnY5�YY5,�8M����C��P�'`�I��0�?�~�����^�2���(Ju��'e�rbd �OD$d�d�T-���H�s���0��Q��g��s�>9W���չ[�j����`K6� ��af���,00s����{��� <���`��IN�,Y9��
-u��r����<���e���./���������{��IҾ�=<��e<w����䀸�}v�v@ �o�3����v��za��w��E���	�"��3�O1����K�?� ��c2j`�!�p8�N�-������/=��OPÌӧ.bu5�f�&����D�����A�~�L��!`�.'~^_ =w�bS9t9�z#����P8,'50���C��4��Ʊ�+�/m����S�8��&�v0"���g�︡��hQo�s&�W�Ҵ����Q�kh��*P����F�4g[v�g�6�ݬG6����v۸�Ps���Obm}E�3��t���V��^��v��>��݀������8pp>����n�P��~��I� �u��Jl�a�D���E��y�b�F�6t���	ٰ�h �kȔ\�����s�o�<��2=��W�ß�"f���`E�2Ma1�{�Ɣ3H~�f���o;�����[��فs�I���W�&�P#;+�����{40u�&����}B����H�8v�#i)���~al���T��/j-�l;0����ќ��L;6uRu����2(�Ij�Z���'5�R�����������_�/���8��Ѓ�51�N�w��P�y�y�~��X m�B�V�&�t�#��te�J�X�-���b0יV�����G{8?��x�����ә�k� +D.��x�ɪ�bb�"��P��0�E���@MNj��)�`}ɫA���5>R�c���"�{bӻ��u������=�".�7�I���8��#������%��a6=��,�Z��\4���ӭ��sd�o��������Ϟ|r������s߼������jx���::����<�T�I��B4�0�m\�/<�Ks3X_�ʫ?Ob���Vø.�\�Sk1����[����#/��\m�����+E�G�4�hUj�ynO>&�z[�*�����+e��KOc���@�����06��;�P0�D,�V��;n;�_��q��.�庶���_~�/��Б1�۷����6����z@��u�L2�+��SO�@��䤦?\�[�N��8���O�B�V�D����X,���\�<'����)M+0��p����-���ć`���#�:�\}4�mM��w󡡘'�����H�/���f�:3�vfID�.Ć���c	IA���f��� pG�ſ6����,�-�(�;	���c������R�?Z�	ǆ�5����r�q��!pE�.d�kop�(��Z�����z;kU"@�ნKV�ty�<m�ݶG�Ė���qr�����a�E� U�ӗ��Z@�o�c�4�"=�Kk�^AOcCQ��9���iD�}Yű)�)F�k��ŕ�%<��I�,�T��C�Ĵ�\Й��ȴ.=��G`��-Z@�I��T��\�]^�~��r+W3���u�#1����`L9 ;0�u� �mK|\��ౢ(Vk8s�2�:}�����-��tX1�׬bl0���7�vZ�l��3�.cfq]�7���#Y-rzi(�b��A,�H*�S���F,�}%{�R���~u���^?�s3Kz��4�A�)�*��Ɔ�طg;vL�(�V+H�L3+A����R���0��C��@���s#��G7��\lH�z�1=G%W�¨Rkb�PW0}�O��E��/��%*?+�!$�p�    IDAT͆@�W�kClH54�|U��d�L��T!Kw�z�Gѭg���[��X4���Jm�����3Q�vᥕc�<�n߂����D�n:� 
Q�����Z/��ř�%Ѽ���iLUk z�C����J;�\�FA���{�kkޞ��d�@�ւ��1.������E̯�s	Ei��C�CD�������f�%��HЇ��al�:�x:�Fx���xaV�%����9�+a�DJ�t[��!h�kBؔ5:���x�7q����!`SI"�P�N�5� �'n
�R3g_��v
�,�A_���Hn�9�E�=��D[�F��G���I�uQfA�ZJ��j}�����r�>Â�_tk�L��_�4>�׵ڰ�D�?�T,�����E���rHz2�{DHv��h��hW���xF����J���vރɉ�����S�L��j��[a�tj3p��d �=��t�_s�HC%�ۧ��X��y��J�M���X�� �{��+�q�����w�����-O#��IĊ������P�R�b|�����{�혞Jh��}Go"/�NK`LG!�N��.c1I��s�C���Kp�S�I6u�v�1�Q�+̉�!�	ʫ"�J!�4:���xF�}'�/�ZJ�ak3x&��?��Ԁ1������Em6�!O>����G������!ٷ�VŅE��\9�:ξ�
�kX��W�hW�
u��H�FB��Q�Bc���}��ͨ^.�Q.�����@kv�wDH���0�O�?ۮ���p�����؈��2�d��FB�<���tI�	E�Ə����\p�H��#22�ԶiDw��Cxkq�<�"�8��V�Ӹ�λE"Z;��G��B�DZ�����n_�~}W-/�{{��Vssw���G��o�x��������S{#��?�kš��@�E�ih���	�C	�p3����U�³^ɨ_;)�/]�5����`bH�"�==���ҵ���KU�÷^ƙ��4����05z�
ʖ�"�mvC@���c�h
;�GQX�����:.�xE�!�C����g�dC�D�ʥ5$�!��}������b��1=o�����㨕˸���|�&ټɝ���imH�P�zI�����*���66"S�;DbwJ>���H!�t"�?R�:��(�#����y.�?���x�Y��	"cHn�)/��P���+�A�a�l"�0"���/n
���=�T�X�p˗/����)�Nd�l�S(O��/��&gq&�*�3�s�����o&�ȶ�c�����~��Ҏ�{ 6���Q|���Ɖ���M6l9:�q،ln G��tNSO9�$��ݫK���-Ca���TxK;+�Zۍ��x��斳h�9�6��F�f�6[z�]ۇ1�#���i��':Pot�����ˋx��re�X��L�d�`&��F~_��'��&�%f�a�֐���D�Y\er�,��7W�+y��j�&Ǳ��c���x���Xoci�.z��Wf�/W%���:����&g�nI�=zxұ :�:���G����WpavA�
���a@}6���Ω$�������Ug$C,��A.-���
R}N��E��E(�Ԕ����v�~��s��߳�i�h3G�L^�LCmt�-50�����e����hv�&U�V�9��d؏�Q�MOP�ܓ�'�28+mTi�:��������欓bh�8e�k(���y��+����'����n�M)��x����~GN�!��k�`���s�y�v�
N_����|p"�>�n�������5:� :=?�W�8q�
^>5�R�����'�����²T)�T���hY�:#���[0=���T3
�^����t\xC���St��pˣb��Dg ݎ�C��L�chh}��kE�__�t�VW�L#���jd (jގ�q��p���P��k1�ǟ?�+�Y�cC�y�Fh4�\��q�q��5Q�>&d�F��nsa�4	N���8wh(Π�A�d�i�~;C�k��Jw�!`q+'�m�k�������L�{�QbgO41<FOf6J�H9�-l::D�A	�k�2�y�)ds�GtRx M>�	#=�RF�J)ò�	u�C�v�L|t�|n�g��i�j�jقF�P���$����1�y-��f�b��q(9B�]����<][�6�,��������g:|&[���38�(���9��x���v�>T��m��n������C�ݍ#��KP]�TЪ�Œ ����ءrBM[_0ͥfҮ�\�tXG���&^c;J�D:�I!kJ���XM��md29Q��ȼs�.�޽Cף'3�>��6¡ F��߀�,��A��S�z�Á.B�����i���~5��k�S0�g�{O<����n����Pb����
UW��<W��0���UTYu:�z���14����B��A-�����F��Ok.��o�usYt�#���Oq~��R./t҇IՒ��X�6�-�'��An�L�G�o�E\[�ZSk��Q�_��LDy�������[�"�SHON"26���R��7���ko����x�g���_G��ħ��Kx���(�=�F���Ā���v��^�Z�����&��w��[���>��M���	T�g����g�z����'�x8K����?�ƽ����MA�DS�dd�i�߆����S:3�P�z���,f��h2�����D�-&h�U��ZƗ�y�g�hb@7L�c�)EŜ
�v���@�݂7�Ŷ�lIE�*dq���p�سX�9��]|��fA��@��^A̤�Ѓ�XZ���Q����z�~��4��fV�E[Q4'^��x��9j^?je�E����ӧ�o}�/_���68p��c�a��#ڐN3|���O6yq�]& ���C�|����?�,�כ�&���I ��@<9�������A�zN*Z�"�R�����1��M̝9��gO��@M W����pP ��n�&�B_��	`�����k���P��?�1_Q�8x0q�ux�?�P,�"T�n�}#��{'�٣��h�9��N�b{�4����C���*]�gC�5�MatdÃIAÞ^M����� ���!��'ܞ Z=�ke,,�Eʗ����Z׃ɔ�ϡD[�bt�"�,OS�x�9ג��enA�J�f�pqv	kk%���=m���z�x0�19>���wb��V}@�ҒƁ��?�Z9��&G���]^s؉H�hĤo�aȋ�Uf���N_�����le�I����x���.RQ�pp7�m�E*7� \��F˫���C��u�ɳ}r�� �=Z�����I#�617&�RL�9�����`����,�Փ�E��Y��A�����Vp7ѪD�ڹ}vMbd(����c&\�I��\�w��p��P7Q攳�E��>�Ncz�(vNcb0��.,T�-��}t���WKu	��Vr(䉦�Thp��|]��^��% �r��ܰ�4�/%ɵr�@o�� n;�.N�˴S�$�Ax!^�]�s��ą�EcI�����Q�d2��n=�]�)��eT��`a艠��cvn�^;�7/�#���V�9�4n)���FE��pc(�R�r������w�q�M�)!V
��ƻ��Z����\�ɳ�(�u��`�;-DCA�S1��-u8G�!�1�N`p0���|��ӧgx�������&�b'�o!���C�qp�V9��+U��-x��]k���g�)�J�*	�G��n�|b;�p�m���V�� �1�Po����wc߱o��v�$�	p�=c-���h��wRm7��&���=�������~�~���c��4J�n�7��D<���4���}�i��Y�~�Ay[t��E��6�P��AD͚����.�PXBmmѨe�,�C�ȅ�ڲ]�((fdk�L�e�A������m~��E���5��ϔ��_+d�tQ稤[��-y�MN�}A$�i���j�dR)�lʤ�Y����GċF�h��� 또衵bYg	�$�$�g����t�ph�I�u6��|�{�R�'v��s�PX��;�T�����1a���t##CI#����_��v���������'��c�=�3o߾=��۱cz�\�?�8.���F��ӻ�qǝw�=q��9d2Y�KU\��E�VŖ-cL&ЪT�_\���<<�&��>�Z��ɠ��(g��V+H�����81>$�x~m��e�YQ�R��RI$�Q�Q��+�g�ٲ�>bXl<��ˣ^%��\7R���w���&S�~� l0��r���Ve�D\%5�b��޶���Y�LF`KDeF��(�5}n)��ky�[-୙E\-V0�g/~�����^Ժ������سX�4P�yP�V�%V�P��R@]���>"4�,e������������?}868t��?���3�a>�����FQ]M�^����΀��o,����)0�k�P�e�T��\�U����n/^=���������*��7҄����{]n�|6e��)�C~�-�
+8��8�Ƌ���ş��1�>'Ђ��Pb!᣺
��;�q�������C�pÑ��y#/���X$d
-{b�iD�\��N�_���믿��~�{�K޶���	��Ƌ��U>X�'�L��1�	.^:1�Z\]Z��/-��g^ų�N�4��!=�ՖO�!�?nh
n7Ztm�[9����F�~M�Zj���`��\>�&�ͨ!ཥ{�l��^�>�l��#�3��J�{0��������Z�X@��w��O�
 ��d��aG$H�n���M����؎�̵�&�rz_��Ά�p���o����mc�|�ۜ��0�"匱)hfL���s�Q�[JÅ�\+��lh����[��2�S[0�"u��b�U��Հ�G��	�aC����	t��8��)h��@�͉�s�Ӆ��J%��3"w�ϗ��S��i	�D��X�R��֟d�A۶�#��ϭ7 ,�v��W$$�0�!/�tJɎ���D�HX�!��XtO��`yh�i����QC�аfe�@V[��_��ª��VH0~~�͑��ST[F$l�W3��h��M\^Z�[�g������LD�i��裎V���4���q��>�t,��DD� ZO��������ui~^�%��R$cH���u�Ɩ�ۖa�Q�2��r�X��q���2f��(0��O.���{���`�f�7V�b�Ԅx�\Ԉ���8�E�ܰ
�^?-�P�V��C��'�r8}�*�:�2�҃H��B㪹$=-�{�a<t�~ԫ*z=_��Wf�����TI���B�6�ۑ#��f��F�"�d<"�F���Pԋw�u��"ȩ0�9��Q����N_�Õ�����^��,ko!�A<yŹ^���H���D���\Z]��W�`-���X(�@����*�%��]�:OO��e�gE�\��m���)/���+�:�V͞[�!�&Ҷ8E��	�r��"�LeM��Ї��i
�}�G�q���_��ۺ��h�ӌ�$�{��蝜�o�{���� 9e��|���ޝ�B`S07^��?e�L��f�0��8
�,^~�%Y�Fcaqۙ���9A�P0�����?�
G��y0�Qk���A�h�`��Y)E�t���u@ɱ����9�O�u)@m���=ƵK�R��{��f� �<��U��d���L�_T�P��k6�D[R��]��i�����ф��H��db�!��-J�}r�e����G���ߩ�P��*cSʟw� ���1br��I��>��q#j�AP��x��Z�� ҵ�]o�����_���|���_}�/T���a<��;�K���J~����~�RQ�mw܊���oK���>�'�|Z{q&W�`V�N����D}&��H������z�/�y��~���	=$�5�_}�6*+k�-]ՠ#�em�p:�8'����Dq�J��j�2�N��D�\A�Rٸf\��R�>pݐ�f�:6�2����y,Fl.�*��+h��#6�T#�aJ4�p2	w$��7�+�".�q~%��L�H�o������=۰���׾���ԋ�t=(�,�Tj���rh�#���Y�a�y�f~��>�����'�w�����'��ԁ���?��@"q讻ߦM��z�^nBl�ItQ'���� �
���$��Pz �N�W3�}�.��y-rf]]%�z��4�hy�8v*���.\m�g�L	~e��9Tp���5�v���������dv(�^%�%�qh��[@�.q�oP�����ӂaC���-�����D�[�p���p���e�N�16:��dRi�T�+y��f�+g�Bh.�)E�/��j��}�~\�����(�,�����0�������|���Ɨ�>.�f��$�M 9�Go��u$t�S(G��b�g�'�*�맩�ϭ�>NK9���j.��P�jg�3�6S`��������m�����96F�AKZ664�Y7aV
�zmxRQ��F��=�Z���w����l��L�K��	!Dȃդ�f�Nt ~����g
�;>��JEל4��;�c�/�5z�W	���Zp�i�Ǣ���69�a��-��XY+`��Uܲ�طk��\W���c��%��ioIj�������)����%��0�l��6}�e�kփ��Us�uQ�����(�L�@<A��{��H�RC���M[_=ģ1]C¥�JK�P+@�M����̕�87��r�I�9!���=�G�H&��twL�3%�@�S���g[]
y��E�b�]��uhW��(�Z��v��F3/�Ͼ�;096��D�<��.�-bna�
� |� �tQbz�b����TZr�aS��ae#)��:��'�6�	���ԑ3S�RG ��@Tk�K
 �Lϔղ	"�P�t�.�����X`�V��l����oB|�wnv�b�%�0�֕v�F���6Q6p�z���F8�g�wO��eH�g���#�k����![i"�Ji��*g��p��}x�}7�R)�֨�����%���v��?�N����m���F��T��mY����ØJ��7ioK��ۥ!��zA��:��.�\����*�u1��Y��#a�¤K@���p\�[ę��X[���F��'04��֩A,̝��oz���F�����Z&�'1���O*��֧��!�A�
I�%�����9��3�yS���Q������	�)6-�]���;�e���4D�6֎��d7�_VS��&�tc�#��L����@���oTJ��H�Q���ꫯ��N���U=�S8�,�N��@9�ux6���b���Q�ca�8]�_D.W��m ���D��B96=ܧX�K{�1�K� [StҕE�2�q�N��r��{�5E���t��vP�Yu�1���Rp�a�K_�Q�@*����DC*��k��>K�a��]dz��k�g�3�rG��P�t�-��)�L��)j��p��!��dd�9��ٷ*n�): QN�k���?���×���_�;�m��A|�#����ӟ�|�_Ԛ����7�!�s�_���x���f��y���r!߿�h!��b<��x$��hq�;�-x:R*��L�RC�c���^��c��$,ҟ�Σ�YA�Z���Ha�f+��h'�n�R)��=���B�B��d����e@��@=�=�j�z���Q6����<Ȧ�B0ArhHZ�e!����,)"XA�X�vG��bǍ��6.�P�������w"0���������K_}�fVPuQ�%"�}���-RBe�n�M��iVμ�mw|���ÿ}�Ǫ!��o<s�>������C����g��`����=��6�Pf߃H,��h�jc�~�}���m�x���a��
n��NL�ڃj��D�N*MX����1�y�u|��Oaf�Wxnz���Fٷ�6/��yhq.N=8��|�I�$3��ma��[���q�� U�-M�h�����%�������?���j
c[�1<���p
{�Mc��-H�⽱�S�+�I�-S&�u�a�z�5|�������;��7�`�mX��P47uN.����6��'��4X    IDATTZ(W��Ǟ���gp�r#<�c�7`xb��c9��
��X��}��-&�Rsa͘���k�أ�����ʅ,�;���f�I��^C�Q�e�)�v<0�va'q7��'0�&8�um���ڦ�=�ƽ�y7�!�4|����
؜Iq_�Zl�w�ɺM`��6�mذճ5LT��j: m��ٜ������@��͇�`d�!��,�C�IwO�:���]�Ut{�Z-+�b��ٙ��/jJ��I뱡!��E��GC���{M<�A���IAy:��(�\XX�ayuM�'�� &@ٿ(��n|xiy��:��ϩU:����qL� �-R-�p��QA�h�������OJJ�RM:���dJ��^�ciPS�\,J���nI�s�v�@*a��]6�nS�(n�B�.Ԥ��u,g
�_\G&_TC�X�	Q"
��秸�S�����7>2���&�J�f��x�Ξ��B8�'/֍�/**���DpP���G
(,H�0>6��-CH����d�n�g�C����
����tx
�u�U���U�E�t�r���ǩ3qu5��7��N�7�Y����gv&�δ���J�f�´�9��ZJ�C�����A�|dF�Ӂ�8�s�gq��<.���"�����γ� ��3���8�~�!�E8E�����Wp��U\],��
ˉ�SNY"�a��R���-Q��D�~9ME"^��:��T��@݀�.�\����f��9������z��^D!�K���30;��z��'����
Z�>�� �I�x�>��X^�E�	���m)Q8N}����X"�/-�����Zn?����p�%��@���8zg�QaB������k��k�nNc���O�^���%;��h�F#a#��k� �k��db�V�|��׆��C51�C��c�'H�B��(J�eC�u�8J�"�?�\!o���4j�>��B��6��\�\}�EQ>ʭ�'�~v�[�m�ԶI�o���ŲN�9Q7<y��d$�@ ��6���B��dêtk�F�^0I�ױ�|Ea�	�s�x�ו�?��Dar�;�l�'p�����m�>s����fq2N:#�1���|���&bFiNb
S�Ƙ��T`~��:�����h�,W��s���Z�����E�UD*��J�v���!��+��:4*i�P̮�C�����������#_{DV�|��r~�~S��������zDZ�R����}>���\�̧�Ǐ���pS�I�VU��#�c�\�>?��I�'�HG��z�f)��ׅ^��z� 7�+�n�h������ j�
k+X[�*w!�p�5��azjB��B�R�rE�/��#��A�׋�*-ݙ��4�����Õ3�[���	��a�щ\DХM�!�@�D�݇;D�ӗ���!G���r����?��]���ƣ�L������b_}�	{��V�
&�7�h�k�e�Yc�b��tZ�YJ�f��{�~�G��{���UC�'�z���٧����u��qT�}UJ����?�Dr&�I��L
L-�e�I�߾�'qh�.��O���9:|7�t�����v��{GѴ�'^Z�_~�	\�zJm��1�������B����4
�YI�`sb�-�+���P �R��9��y,�K	�^R��E���⮹i�c,4B:��ō�E��Ci$RQ'059������G02�@�]f��"u��F<`n��]8�8z��޳S�~���sgRc��B7T×��A�_;�?����ﾈ��^����SX��Piӥ)��,���/�M�t����&0��Jh�藩{������Ϡ8;��zP�0��ף�6U0,�9qv@(�Y	��&��ZC`����٥�u���;[����<D_4���jL3p�!��p?g�ƢcA�����h�bY�1�����D�|(��,���EG�@79(���g�ɮ
꥾�ORAX���nB1�-R �r�,�j:Rq���<jx~��O�A�TR�p?�K%mb�r����=�g!&������ghQ�I�:m;q��A�%È�L�'T>+&`��2�9c��'<�+U�|�es(U�H���ġk�6nN����i��&��`�t2�F��:q�>D�1��1��b���]͉�_op��7<��_p�iA��p��FØ���萊h'�:�����[Q�Q�{��5L��:t�`�g� C��~K�
x�X®�ea�	�I�Ɔ���8�˩�@���.\ҫ�E��fQ��� �Ei*������|��A��M��Xtj!T��LC���gq�ڔ���p7^��'R���^�3%�y�D�ي+�RO�?�h��,��16ǭ�^�T�..,��(�8u�<�\YB�B���\�L1y�z�9)��:��w߾HDج呈�1��b(`Ic�s�U���x.W�*$t�����r�����<2�ZI�,n|�F�!������
�z�����o�#=91��w�+�V��i5�s�U�Z3D}��P�UW�֔��7��4��L�,ę_D&�Y%2dx"�lr��^dL���iL��â��Ź��q����Z8E���� ��Ҵ+!��6��ͦ�*;��S�;(���M�a��|]5�N�gGtFx]��݅����g�U�Z�s���EMq��H�(ѭ7E�3	�&o��e��Bj0.�7�˗/��P�0��nCNF�줍y��*�;J��--�I��i�p3.�.�5����I����z8��#�/���
`�z	I�١bB8��^Ϥ�6�H�����.6l�ȳo�yZ��~t[]9�M��_�Qw(�L�)�.Rgi�KD����lv�D]x��SC�� ��Pc��YB�,B�y
��w5��(��p�������m�x�|�S��׿�u�c<�n��V|����(C���G���R}����w�w~��5t���k����WDVI�k)�Y
���m��X���H�����tЏ0�z-�uk��'�k�5�rںe�۶b � y�H��
��<��>/&G��$��QN'9�'p������W�S�T6�=���?�=�I-��C Zw0��
G��3�{d;�P\v�j0��pG��R��@�l�ky�Ã�>����!�c5ˍ���x��sx�/���%d+��J;��
�P��n��e`M���1<��{��_��_��B��������|��j�����$\ͺ�Xg�8�l.j�����0ȉԶQ|�����x�����k���u���{PkU�jW�e")_+���{~���R
":8-�C�f
M.�_����X�p.v��,9ODC�3X��@iu/?�.�A�Yj%mJdC�!�i�0���Z�ŉ��<��z4 T��p:���Sسs+F����4��)5S�z�����(泘ޱL:4�M����4��+�9��:�%GvN]�����{x���HN�ǎ�c��ë�/��"�L�Y� �1K���(q��b�K���8�Ǵ���+X=w��EX�ڍ��T>�?ѡ�O�k�7wX��.C܊�!�x�Lk�UCJ�����)��=t�Q��އ����[W���Z�3��1�99͞�{�J�����_�4���}l���7'�6��"̞�qs�&�k�099��"�� �]��`�
i�Oz�H���V�XK�]ȞF�ӱ�#	��yH%+�~�F�h����z��f۫D_�!Y��;� �5[X̓Q0�)�X�󳓊�1�L���DCj��[(R�Ԑ�Z~5[h�rexش�5���;B,M�!�.�?�#�`��?/Ұ�$���������Xi [�
�eȕ,Y�$k6�r�Ն�괴��[b1�R�7�$��2(���ax=!�xh+,�e�}�:�d%~1�9�o�ը�ݬ!��ar��G�h�5��Z�x͖[�j�Y:q��M9Da���X[����s��]P�����Q;���r
5�n���Y�*$m����.7�6יT�:�e���Ά �a��V��1�T�6����N�>���"���珙�/��9u�6d���ƽ{����� �	�_(��c�c~n>?Ù"�B�Y��Ec��^$��_(�š��e��DZ��LqN��6|�9A�됷��!V��y�zq�T�A�������-9й��s�?��W�"�+#�i�P��v��\���55 �ǣ�=�`i���j4�.P(����K������U�/��3��*)ņ�Z����j�ۚSp;�}�����A��懄�P�":��:���%���k���i,d�n�r�W���5v���KT��y��%ҧ��&��Ҥ�SuN�����L%�X����o���ـ��0�Hi6��4ѭ��rPǜ���`��֤��`:�b�{H���(�'�+l����}*:�ϭ�r�g�9�����ý7��D��Z���/��iL���%|]f!)��E$��?��<���S��b(ML�&EZ�F��	�κ�д[�j Hg<f�,�iT���Z6�>B��&�<w��xF�y�k�?΀66���n6�.DU�^9�l�{5<K�/,�����Q��h5����=��G>����.�O��|�ߐ<��;�����ɿ�k<�oJ����S��)���>�` ������G5L�~W�+hZ�*e�x�]X�2nR� B�3�j��+%Q�9���h��5�[��� vL�a"�Bq}�|���C�RA�U�����b@a2?���Btz*�Ir�7�ܢN��L���-�\P�H�_}�(i���<l���:3�z7�.DFR������7�^����"4�C; �}��A,�w��{O=�㯟Ʃ���Zh��@���VWNFހAvi���m�iHf^C�������?����7_8�����UC0:��lt*a0����9�7�_��C�ڐ�w<a��q�ﾻq����t�
�|�$Fp���h������4�#���A���s�/�ӟWs�c��@WaE�_-�"�g+m"]mi�o���aaі�?�U�s���S���^x�;�@;RZ�lЯ��]�+	��Z@�v�jI��T:�P��!mq�#A�~����)LOOcr|�x�v�F�c�<��K��1�=�v�J�W�:7lt��Wѵ)KWM��<�Z��ssx��E�b(��87��\����	u�m�RTı�����! _�'-�(p���V^�`���s�p���6*�V=�)���'�f�jN�lm�G�' �0��@��VZ��攚��ǃ�������$����hr��ٱ�sH�.�G�?�BK�l�|���@�Y�kA���<�,i���^+��ÇɎ<pk�q��$
�(M?�czd�L�9i�磆�O{��i�	�D�wP��&� ���H�N�rS����J�Ɛ�
v�=i�Y=I�g��������!���H���ÐT8�{��m�<*�ɝ��1�J�}�sIZ�2�Ic���z��#U����S�C�HK��ɍ�g!��m�R��Zk*������,$䳭��N3h uD�����ę�v[6?���~Q�������sȠ t"��6jբ�nʵ͵��M�I<����1Fl�}���bmmM�|��=����%Z����QL���*������=�u�ϝ��\�����m���j);��u�mNa�����^]\��jmX�4��}��I�6��%TjY�A:| {voמt��
��t�L�� �~>�"+_;��r}�>�64:��� ��.��aj< �TK���
;��h���0BK~�`8�h� .��ȬgU��v0FZ!�) .^�ًW�J�^ϭ��&������ۄ���`�L���'��f�\��م�[}DÈ![�`~iU�qf|N��������T�������_,86ڛ~�>�9����w��ym�b��(�|��E�JT�?ژ8M�66LZu�.���i��7͉��$?�<mj�$�1�2�j����l4��<\�n��i7ѪT��G]��{����GMa�;wMa��	Y���&�� ��L����C�����÷w�!����.
WWHQ"GG��D����?;;��0�/����������n؋J�����5��64�Ȑ�x<�}����u��z�ͬ���u���%��:Zg��셹�=�"��E�P]��&��_y��#�NP�D�23#�d<�l&��Z�h�z]d���u�1�|14�h�_C�����A��/���Ͼ���N^���>*g"�N�Ft�=wȁ��O<��'O����&�s�=ǳ/��/��/���+rW�!C�� K?�!A�s�h�Ҭ#�c8J�Џ�4��Х�F�uN����hM*��2Q}A"�ԔQG����i��YGne�b�3DlD"յO2���3�P쮍��CP5�t�j�^�2MAzpY^�,�jZڌF	�q�{md�%�[}�b)D�	x�f�j�j�6�k
ض�����L(��@��:��}�1��-c=WG�� VXa�e&۳q�]4�o�Ԍ����<O5��O��=�~䋿���6�����!������-�����I�U�qJ�B�Dg-$�.[SD��
".�RCp�mסWf/.��+bppP~���ʷ,��������<�����R���d�9�1^�t�PC���5.j��.$?y����vTK����o��μv�䟐���M�pʊ�1�|����A������+QgW��*�r�������j�}�y�hB�� �i!`��1�r��߷S�Ҟ6�.\�>z>n
$Pз%(KJ6�/=r
o�[F��B���|���]����ot@������x��G��-ѓ�<fO����3�W�J�U����D�����3�(ͦ�( R�@��Ŭ��m6��x����N�q��[���LCpumm;Q�PH���֕s����-Z��>�γb�w��2@�4����s`���Np�������;�~�<p|�up�!���vp�sTh�9超����j����M��c/�i<�~�k�g�O!3����r�����]�E�3&>��Ιr���+:m��o��^�𾈊d�٩S :����4�g��Si����>qܔ6ayiK�-�¼W��#Wӆ�IQ���^ۮh�a���''��s6��S�}pȔp���ҫp�.�~�>�5>�@�S+Q-LpC�14f���2�ev�#��d^����$��pLa5�>��sr�Ϧ炰�M%�L��(��a�E��d6��2�ʙ�I�1�6��gC�f���Z�EoǬQQ%xo�A5_D)(��ǵ�9j`Zuԫyt{5���a�]\�<��匚�h4�)8���7���/:��R9�=�{��P�����m�(�汴�h(!���䗅$���59�޴_�ǒ(W+������&�&0�e�XTڎ��%�/-I�BZ�2������M7�M7�0i�Bz�RD�Ҡ� �Á��"2�%,�籴�A�ц7��Y��|M�x����8�2ǭD��Xn>��P���恄s�9���%��I���{�f'#���}�F�4t��Wg_s�x���GyM�;S#V5��� 3�U�T���a���d��U����J����S�cmyA�d�P�J�,���EL&���f�T�DD|��_����.��'�!��v���WHI%e�L����I�醳���m���8�;��u����Kp�u���h(�͘vB~\�]�?}����w�@��B<9�ip��������k�ݦC��0�އ��y+n��0҉�PG��y}B�1�G����q#b��ba��l���q�"�9Tkh3���&%@����C��k�����cnv	1�������f�k�~�w~�x�v��$71��^X!&����3j'�X1h6�o��c���~'N��/���B�n��x���B�`���Ǎ�?��P �mC��s���X\�}��s�B���<ڭ��YXC<�G��G:5�~��e�W�U'9} #7a�D�6ٌ�A��o3 ݠ�fXi�Y��Z�<�15�'<+��{-,�����#�Jcxh��4��0���k�B4�s7Fv�C/1�~j��'/���'�ǋ�^C��W>M��4������8~^b��    IDATc�ϳ�::j�H�%�F��n�����}�����b��?|��hC𧏼|������\����D�\L
�x�:�b�9}�t�� �e;ǒx�����[�����&��qs)ReC@�;k:��{�|�����<�1�^�`1�ž��=�Q�ȀN'�DP�h��T.��_��=I`��l�N��^����x�<@>�Bi��7�^ZŸ(��aE#r�`S�~�D!=�;6�g�m�Fd`09NS��v�Ѩ�U�#��!7؉����m�8��m�M ��S21))���_^x=��}������/O ��@$�/L4�"d/�L��H�.�X�x,�>YBa���+�"�AHn4�%5s�O�_b07%�z�&u�T*�S���̦�>��l�ٜw<�ʙ� ��)Z~5�NDq�=�n ��! ��1/b᭿��&�׏6�D�ݙ@r3 ��M���I��D��{x�8S�%S�U؉�>Ŀg5`0�s�"j��|��ۈ	?�C���M"v�F$��B���(�א<YM#Y �I�lN6Q8�g��i��i��-CVv���E�f\rM�5uDߢ���tz���g�n��|s�ߘ|k
Kʘ�۫�н67l�0n��7!���h�,)�j�fN�g���?C�Y���<�w5|��Y(̣SQM�"S����tS��1'Eͦ�M�mG��޿YC����Zu�T:<r�?���hj���ϝ�RO���b(�{����I���c�G�'�����9lN�7ܖ��6( )�>e��ى�3N��IPI���3
)�.�y�>��j�|Q�@8���
TsWl;a)���z<Ba���2� ��-"���Y�X"�����T������R;ʵ��e~NR��=�J��6@T8�z���EMȎ�#�#�vU����a!9�֧N�ѳǴ��z^�^�# @��a���@�n$���}���ZW�\��ᗹ�5�Ú-��|
o�8"X���cCp�b�������&R��.d���zQڌ8?���k;T$�z�<�����i6$�Vrﵟ�P��`:���%�%Q��DH?\[*0�Jb����8w�
�
�t�
�P��Ѩ�p��C��G~����q�S�)��ك؀�i�glz��G�٤b��[4����C�<;�?�=�h�I��@���M�����|/��=�U<^���h�FE�/�>�3?����6�xx?�4/�QN'��d��p���&�kC%�?�����h�**�a<�3wXg��h��d �>��0���|�<�«�-�Q)1p���e�p� ���;����M>�	�8�\Y5J��Z��h�<��H��-lm�@4:����Q<�w_�Z��V
ylsߕً�fY��[��!\�k'RJ+�M&�k��Ye֖q��9d�W�����߇X ��dt
dmZ�SP\D�hJ��Z&HJ"�U04�D:!��YeQ6M��m�}S��A��Q�;�d6\=d����ʨFrx�d�XWV:�����jǅ�zg�p��9�~�<��`���� ._�f����|?ls�V�\��q�SD��x�}������?�yo�����hC���|�����|�Գ��F��$�	!w.sj)Y��m��qc�� ~�����Ƅ�_ZE�TV��S�@���+���s����(C�����'�#���h�tKv}�ЍK��K�	�7����H-b� ���x�]B,�C<�Bu}�?�$.�8�Zf���[���DI~���#M�b=�G4G<�ւc'JGA�#L��G/f#��D������`*r(k��r�!<�нؿo���1Ӆ���Vn���ᱧO��L�kMdJ.�"i$��55�D���ϵ���ߚ00M�'{t� /�Ԑ���)��,������.��KJ-a��������"��7����z����Hx�X��DRrM{�hC�XG��Fܘ__Cop;g�Psl�"Ûw�h�@s��7�y��s eN�w�h5�9h��F�V�o��Й�I�����Z�qMɩ�\�!�k���j�ɟ	�Ѽ�1�[t.1��-����o��D�v{FwD��Ԑ��i4TH'|.���257.1*�mk\��P�VE���F����'즀�
�k9��UG���p�L����.5�j���b�)���6�L���kſsP����E����P+�i���0���-j�B�LPfo��ȧ�ܦ����x�w�9EU�a6���R�d&Nא�����;�J�MɰΔ֡��&��R�)��arl'9Ø���Fw�v��㇛6���f�#'�_j,l���)״g��� �i"�$�e�X9���O�<݂��e��Ws�k�� �:�:h4���Xt�"�ד�����4Xκ�wS�K�g��Q�LU8���c�;D��Ա�`A�$A^O�Z��%��ѱI�ܹ[� \���8`��zx�D�4�r������A�[���;q��.]�7޸��.���ĵh�k��c�s-c@͍��4�,W���#^c�\\[7��b	T�R�0�4���ݔ����+�cf��5���h8�����?҂�#'�������_x�\�@ >6�ժ&�a��vlZ�0k�=gl:m���q��7���p���R�F}����6�M��m�A����}S&��D�m�E��K�ى���l"�+�z���!=�l��/}�[���:2��\{>�N���}��	m!��<ʥ,��/����ߏC���̊�.��z����{��O����)\�~��^'C���W>�.���lL�-��7-��4��R�������7é7����+]��#��W~���mo�Ig:,����:�H���<��������U�����ￌ�����y�d������=t9جЭ��jԐp��}x[�i4�9�l���I%cj
.�?���3r,#e�Oξ�':P���«i �P�'�d�k��tl��yr�����e������j��:���¹�^E�>T'���bhp�X�h�tV"+�!2:
w:�\ߥ`���\��󗰚)�W����j�Z�IC=�Oȸ�1�X�D��e�`��j(h�t7_��}w�S��K��&`����6��/����ߖz�����}3Y���%�2��D�.m0���*a��m#I�����ۑ_X��S�0O�ྜྷ�E�]e�7�<`7�������/�Ņ&ڞt=t���&2S"v�|�X>u���-3���Ð�>��<�u���X�.< �y�+%��Vp�Q^�L�,��S�k[Z���WZ��P����h�RIŊ(Mz^w	��b�DtM�p�H�aNB���C�Q@,������wb���������ե&.\Y��/��ϣ܊�o%a��Ix*ΫF*���=s�ІO�;7Szޓ�ۍ%��k�~�Ds+X�0���˨/�ʩ)#�0��R)g�������3�s67z�sj �<hh���K�4Rg�poj:>7泫h�<zP��Ξ�+s��7��fm ��YC�����#T�cy�b�<M���tж����Lµnl�9�Y|sh�����ms5̤���G)���iI ͢�43��j��6	S�f�(	�	�S\pZ��:�	C�Ź� ��g��5�5Ź�*~�`hk1t�i�j>�S�N�É?�]�l�����7L����s;���r*��ڻm�Cw�N�vҚ����;M�S\���,' S0�гiT�S�fϦ|yY(����~2u���6į����_ܾ�<�L���k��L�c�nNa�8�8��:D� =\lE6e<08hq4.
3�ٶ�,1h�,q%�p4�hV�ۙ۸D��i4ύy?���bR�I�`�_6��Nb[.r!M�˺���FM�V6��>�咬�����(�^���@�/l<6:"Tz�$��B����8�LZ+,��d�ZZ¶�T�9�a�?s�e�}]����4� ؛XDR{�DQ"EQ�-�O���l�qދ^b-/�8~�q�$�K,YT�Z$�E�I��@t0 �o����������<-��Y�̝{�����>��w:�D2��K`͚u�Ӈ�ʒ�gP�6�L��/�u޿�T�ꠇ*VOM��K.��T{������Q���i��+�f�hVx�<�zO4 �����:t�L�6�s���W��Y��`s�@l{��#�L�^���p*Ӡ*y�D�GI�!傒ƹB�׮V���'Cu~��t*k(fݽ^�#��2�����eT��p�-���~��᪫.Qv�Z�NZ�)�	�2��1�e5&�8�Rɽ�R�ܿ9ߵ)*��Vș���O|`�hʬ��!	����w�����������Q�cT���>'g[V�c�,.��+^��~�}�����Bł'�:�h��,9-@�:�;�*���(7?x�!��9O�'~eI-��� ��Ro�?|�{�ع}�Dˋ�J�G��k���w�"���F�S��g���$'x&pX���##�3�SK��K���>�:,sG:�sQ�I�d����"��&R�l51�L�3�۩S����0Y���-�cu1���c�?z
I�bK�vJ��RX:vL���N��J0���s٬��t~��h�.�II~4Z��5�{�*���b^���(���L��126�3�<GeLR��8V�!51��-�a|��.��ܞ�x��,�Ul�;-����*I�֛m5犣��Tbs2���3�BZ�,���a@��5���7}��?z������~��W��?��?o�F�/�یr�E�	�����j�Ь�D*F�D��֏0�N�>7/����]���}��݆����t�5N�p`��/k^zmˍ�Nb��I���j.\�) q�]t�-�si�Y�c�9}�;$�˥%,/�����߲n��w��<��xs��[�R2���T��[)�/ 72���ˌ>m�{NXnd�pHSbS $�E��@�e��eՊ#Y�s����w�k֌�*i{�/��_ū{��|�u*�!S\$hD�E<fTWwI�C=�Wv��2F�:X�I�p,d��d:���
J��K��^���νX:2�����+��Sw��ryI%|>v��ؚ��{��O�B���agƝ�$�d���?>����
׿�6�i,2��h�j�x<04�B��Z¢bDx��z�CMf,���Ohf�Z�{#����vp�l���\>�x�����~ ��m���|�������р�KM�ZHIS0��d�E)3qS&��:� G\���C��q^����^�[�#��2�*z��sɵ�*�^�f�����+>s��A���!�McCr©�Ōs�4�GOz�oo�t�st<Np�V������:�I�avЛf�lЇC�4(~��h�+�Rx���FIX(�����܊����AU��^��4�a�`�5�Gz08Ol���޶�	��{s0�U8� c��ϟb�H*�g�Ǫ �'��h6N7�A�{I�#fr�3�+LRP1�z;.��;��k�.���e�y����5Z�Hؾ#3���,c���ۺn��P�D4Z,j��h,��k����,C�\>4|���S�6�"��̑#GP)W퉽>���''T��&Q=����*��[bÂG���K�f�{x���iY;S�� ��_���u�Iq%B�Y��b��	J�Ze�2Iyw��N`�Gu�L�h�G�)��r	I�Al��t��_RB�^�M7]�_�ŏIΙ���l`v����߰w*Ẉ'E���):������mdh�HF�+��c��W�AF�%E���~��n�~�\bro��Q|�����|Dҳ��6�8>i ���lZ�����(���,^w�9x�o��/�9�y��a���0弑f��W���x&�Y�G�c�"���P/ӛ��)d"����.&G�'���A���\���<�8>�ůa����Y	��I]�j�m\�vR	��ʲ�Xm���S�O���C�-Fֆ��◑����i��G���<I���T!`���"�*f��X��>+�&�EQ���D]^F�R¦U�p�i�o�Q^�W�p�6����=Y1lw��T�a�R���E���Zd����ϣ��z��RI�g?��"���0�U��
��#EU8ټ�錳�.�Ig��l���"91�5睅v����"v9��z{�b��<��Q�(z@�,V�y�3��j$�+����3##�.R��f�L2�c�%�z�8FR�g��;~�|���hd��ݟj��?~㉫�3��%��ݰM�7t3X��<��l��Zm"֮�[YF���vW�w>>���5���F�"7X_4,��	�����.>�����9�Zĳ�Z�#��F�{�q���q���=Yrǻ@��B�N:�n
�&���eeF�i�f3X75!��~��g�p|z���K'��S[^��'%�W|>R`x�$�Q��2����3�s�Z'.��4T��S�^A�^�E�_����7n��ޱc�8H��gFO��է33���h,oʕr�2�7�K=��$�<7�LJ�9v�+��*���mT�e4��X:8������2tk�����p��^�2�q�18r�����D��Ӕ�m�[=�+n�VA'��������eR�H��QMf#HN�NS���
b�H��xpC�Ö��4c*5G�G���ɗZ�T@(41��g��4���Nм&���\y�(������Ɍ�"rMʠ�0�3ޤ1�@E������$$z,�JQǵ�{J4(����P ���.�f9aK�����D�wݣl0`Q��d��E'eXD3�a�.F]���b �2�r�M���D�-��*c�kI���A���=��qg��R��>��e@+ȥjZX �4%�b�P��^	���xt�\
��g�nܾ��
��<K:�ty�5�Ɔ����K�\��y�yo�5���Zp� N�fLiSֲ th���aŘ���C�@s�W�3�~�tٗ�?t��3u��G��Qw�(L�>:�L	����5r*�d�W�(�y��Z�FG�����ʞa��oJƚ��{��{�����&:�S�z���@���[\���*?�+=^��*�������,{�u�6���粞�'.\�4�%�2����u�6��������@�۪qe�llԗ��Oca��49͓f��N����U
sؤ�\�^:WЪ�p�W��~���K57���-�~�o���/*+�yE�+s0���~<��>���,k��HqN0��g�=>A���)�%��5'?2����#ǰm��9xTՁ���D�0�R��D�ɛg2�F��&��F�Y\t�Y8��3�\���P���y�0��elJE�{eɟ�'���O��Z�RG�TU�y�Tv�gp����3�2�r&�R���<���s_���#!�W&4�6��*j�E%Q)��UT(u�!Hn��5����3�A`/e�R��}���E���9��Yc�]�9ߪ�8��C���F��n���#yd)�@��n�J=���C�X�R��H�u��K��]�uN.�	�/�M��bE�%d��r���b?A�Mڭ�����-r'׭Q� ��F���踒Ӊ�1��I,��8Z)�G��~;��2��FV��Kcvn�rMU�|��&�@����կ@�Ca���*;4#U:�X��W����g���7}��?q�s'm�?�~�����������?_i'�/n:=���}���w�pZY/�O��֞d��N��~���X�_v)��N\~�Z�V�4W����}�L����E|��cǁ
j�1$����Ry���X"E�R�d�JH��~�b�\`�=������Z֩�h�Zg�e�Xb��i�)]���֮�S*ce�N�?��ݻp|�>�F5ₛj	����5�X:J��W�@eJ@�t#n����v�ȌOb�gb��3��\��̔C:7�~��X	�0ӓN2m��*J�%F�l**:��L�/������ټm�q�1Kj�q��3�W�X9>�:�ҩ�2o��T1AGN�,�G��YbL���1�8����e���F�AWz����Utpp���Jj���%���t�m��7    IDATӤp�Ų{;zD2�^) =����OV�5"?���a4�MƲ��"9 ��{��$�πJ"���� �|�6f���2���v�@A�����H�;n*>�-���$c5

`L��><�L�ga�gȲ(����";�E������^|R-�l4P�&UЂS7��5Ǒ/Xf�i6����2������e��^j��?�E�4�v���v-#��e~ך��q� <�z�9�3�=(�2v����)���Ѓ E&5�M�Zs6��U��Ï�z <�$��Ж9����>��;�����.5� $@ۿ�z�ϝ0�{ʚ9����(T����k\dV�����5h��g�Ϝs�Ϝ��}�᜗�":�U������c���ps���]�Ic�~b=ދd��x��k�גyҰA� �~!T��ך?��9W�5;2��^�A�����υτc�����U���< �@x�w�5E2��x�bM�� MP�#,�h�&�4�N�M���ʶ�
�,,E��_��(���r���r~�@ݩ�K���2������	�@�lQ܀�#���=��w�?	%�������D�=�6�|�>/���&�TI�#_�����I
t��UVy�ڵ�D^X*aa�&��5p�����h�%��*0K�<�# �~�f�,VD�
՚�C����s�f����F=�(�>�3 �Z����܊)�ߪ1	G*��X��U�������{~l���w�xt�V��/|Ͽ���6&�+E���̪�H�|H�b���@���S	��1��k����Ϭ�ɢ�J����� �"��$��R�d?JW��
hXY*$c�0:"vu�&3)L�3�p��r�'b��Uj��3�2���T�SP�B*Р���qV�E���]z���� �ϩa���i[N�i��hn�9�c+%�,����Y��x����q	�<�������j�㨗[��9�>�:�khI>)�Q��F+�G��=Iբ�r榐IeP(d�j�@�S~杷_��>�sχ��'����7��������R;y�������0+cRB'�fr�S���:�XU��b���sq�o�EgN�U[F2�����q6g���G��Q���r��$z��� �&s��i��+��R�綍D>�V��z�j&\ɔI��%-j3�48����JiY��ѱ���($�X��a��:�Kx����ٷW�
sǎ�SZ6��h�Y)R$�9�X���0J��*n(�HԘ���Mظy2�Q��^�.�L�J�����E��B����}�����e=�hfe1d��$�J��	͊��jXN'g�Mz�r��4-�dmnz۞xG�����qU������Զ��DeȖz5�����%�hi�#�EUz��A�Qܸ���&\��۰�i`ϱ�heR �΍�{/��9f��ݬ,�0 ��e��xx��3m(l>��ឭ@
R�j��2��5vZ�س|�T�,x���(�?��`;�f�C�����@SP��x q�M���mt���@Nk �V#�=�;��J�ˋY**]*tp��W��V/4�9��ʹ�ENYp,ץ��W'|��5:�@�8�b,=���T43:�%Cω��"{V��!��~dc�Xʳg'���c��QT���Sdb���VC#+5�������"�5�%�	�D��3sE�Hc2��I�@Ф�B�u��l�(h�'�����)�f� ��i�e=g�Ư�
�*�<�~�M���eߊSc�|�(�=T�Bv�b&j8$���=��*�%UHsP�t=���f8ۡW�`�`�@UTCW+�>�gP��P@kn��+�x�
�,���w%�����m"�f`ߛ�*b����h"�i%��'��J���^�h�
M����耒�&zV�,�
A7�==+�gw��������2�d�P�Ut�T|91=��܂�űv�$����S��UE�S��7���K�UW^j ��ƾ��[����3/��l�fzt���0�)^'�g7�A�ߑ� ���cC��q�E��$rycxe��a�Z�۰^��r����T	�{1��cX�z��`N?��Ξҋ����ŪS\ �^cƹ!uD�i���i�8�J�~EU��UQ��GưR)�Y�Yi)�� 3�F
� �S=T�J�(�ܴ��x��L���n���>�.��O�:�L�j^iv�ǟ����ں�NRtY���*En�6�X�Ғ���W�[�,F��:m1JՊ�a��I=X!pW -��Ћ�)�<U�xN3QK�.ǫ�kJ��j�m1�Mc�1L
(�ۘȦp��5�85�$nu��X���B�j��ET��~��q,P��INJ��4ִ��{�\'�s�R��ʓV��}rM��i�3�w׮[��u�P�7��(�/a��1̔�HM�F~j����C#�Ś��R��}�d�jS���� -;��I�bB'�}�O;I˓�~��ݩ�V�G>�|�]o�����c���G�������������̟1q�Yht�J(Cڤ�S6�z���{)�G��Z=L$Ӹ��;n�y�&�o-#k#��]zZ*16�ā�>���ڋ����:�LW,!�	>l��\i(��S�J��J+���5��nM�Ծ�!C5�BZY�z��T��M�3S�����<���<\�e�$��)�о���SO���=�4�.�/�R*���j�5�p���(1���*����U�^��ι��4斀ٹ
L�����Pr�%R��L��h�pMsB�%�&�덂���r[l���C&���e8�l�^�����K��x�����]譜��͌���P���=א-7g���I��Д:��3-�&�;W~���3 ��M��ͷa�����Chgɷ�˚��1 ��Zڱ���7nj�iOW�	 �A�Ξ���(0�� �{So�-k$�	&fEl& `p-
����X�jieſ,���Y6��>�$�w'ne�)�+�����Y�2�D99�m�=:Pj�7��L2�1J����\���y��a����yp�\sn8�&�=s��&
�4/�3���4�a��[�p�,��7����蜉fs}�x *p'��Y�25$uP�
�z��V�������7&dB��� �^D��k�'��t$��u'������k�੒�5(N��*6���'�qSf��$��Mt�! �;u��ż<��t
9���H1���?��c��!���Bo�?	0�I��H:u'\u��%������C�?9��x��'�ao���uƤj= pRu#4���0�s�Nʈ�C���
MN����W0��`�-���x��X�X�J��i0g��֗A�sO�@�M��H�����bi��؈�g��F�%���gqp�n4���o���0��{/��
:͊T��r�����]x��0��>��K�7���4֬;�ݥ[���3;����q����<� >+�֯_���U���eq2Y�V˘�[�d:�G�C�R��F䍠�o�kT�bZ�ۄ5\�Y��f�I�n&0::�
m�^{����Ie����j�b�@�H���P��FM�ɞzE������z���&��
A�����t3���6m� U-k|g���7������̂X�]�R5ʨ��6*��Y�4i��\A��쑡�K�Mz�)����%m�oԱ��s��+���PO�W�������t�s�RF>C��b��Rq��}��a.��|��i�ԬJ���lUj���>��j��6f��2��b�8v*	A�4�驊EU��kg*^vo�W� ��x�t���J an�T�k3GQC
�USHQ)��Z68oX/ED�w���R	ե%�L�r|H5d_U��Ud�����N�J�Id�	l��ј����֟�?�;�{�?���ӟ����������
�7��߂*Cxq�-*Zq�6Rb�!�ٶ'a�R�R����*�w�M8k]��
���3�,�р����/e��,/l@vtR`Cґ������y��b�NҲ�A��	Ө"��j>�2�H�hqQg��h���C��fe�^�L���L�q��I�}7;`~vIe,Vfh���*ڤ�v*U �1ڭ�d��$�����S��@���J����B�T^��Z��T����d��lyp�%������Nl�"��`�)n[���<�H��uQ���h��0��n���
��GE�2�L[��(p�3L7j�r��ɔ!r����l��,�fzhƖ]�W�~+nx��(u��ulʡ�䯪H��w	:H�a�d��A}�:��v��YW��t��0x��Pu�L$�.Ff6�l�[�Z����n8h����E�����_ `@G	}=<$Y������ �v�l�����/ dȃ���E�"��iX���R`43SR��_&_�Sde�g`f8��)gN�ч��Tq�X�U^<{-��S�^���@b�K�?d���$x���g��CҬ����PAhҶ��A�A������@5;�0ʨ�<� �
թ*}�Y���T��:$@�QQ�Ɛ�&�o  ׽pG�>�Hf$-X�n�lB�+r�b)f�$�hN�J�!e�c���|o�\��v&df�>e4^��h��@E^W��jM�������1�Ɛ@{,�$p�~,���{ (qܡ�fB�?:�ˀ0f �e��6�9n�r�������_�|sJ��'��G3�>w5����/��CN����(p��s:��y�� �jT]V�8��V3��;bjbeB�����~��fm�^O�-�kaϮ��k�NL�[�[��O?��݃�KKK�?4������'���o3,K8����mw�	�x������D����[�_�q��,��QbYuaO�V�ʈ�m��2�+d~61�J�F�Z�
�揋D0\���9�K	��yy�Yg��.PUb߾�8zlN� ��"4�LJ�6�dU����s��(	��Ϟ��D�� ��Q�����H�d�;)Rs�����)9��d�0�B�
7���b�~�u��O�slܰ
4%_iv�Ҿ=�����Cx���p(P(%�&i)�;:�e�cb�����^�4 ^�S��b�}�z>��C�6�_<�H|	��Mn�L���F�L$PV�> ���?�vkFGq�y��+^/%DVV�PZX��	A�g"���q%�Yɨ�k��}���d�Z3d��T!e���lު?T;cS|�b�VAf��x���F]<Ɠ8tb���QdWM"�z5��+I�Q%~d�k����
ZՊ�S��[�(!�(��t}�����(ɝ��ۦ�UF�q�Ve�|�[�����G���O* ��?��=���_��~a��������7����@���+�+���q�v�Mt*u��Ҹ���p�m7�u#��K���R�aV��g�W;�W^;����s�5͞��
D���أh��ή&{�,(۹ɫ���O��I���"B���]��p�Z��%��c #�H�\ZU{�q���� ��P�ʕ�]��&&УT_�I�V�r��5�r4�T���F�d�M �����<M~?��R�^��:ԣMۆ�d�[Щ���-��(��N{fK����&u�A>`�dZY���B�WA�F�	��j��H$i3:��X���{��6T���o�8:�Mdyi�z�Hd��0�^����4uӖs;�إ2����V�kp�����܎r��׎B���J�����L<�S�ԕ��#¹��ȳ�C}w�Qn�oZ�(4�&�����R+�I�4����D�?�BU؜H�(4�w�P�����>�ܘ)��@���N�t�?�q��*8pl�j�6�!ޗ@����*�]KI �=*�|8F��Ź�'����fH���'���9����Y��̜���w��4T^P��=(�=�{�oe��+e���`�4�;��h �
Q�Ș�����Z�7r.,P�%���S�-ЋɝX��@{���~ŋ��J�{���k�3ն*�2��5z���ԃ2z��
�T�B��ԦT9
���r�r6(4��h�$��x(`�qt*ؓ��ҟl�7J�St��T�"�ۘsx?\�*���RA�#�"߿�+�R]ܚ�ɵ�����!�p{O�<���d �zBk,TD7���7��� yH�1řA�R��<��������ak�j�
��SQY1�R�_	��%���ʔ&��� E��
��.֏0�I`����S��x�ݷ����ѹY�x
�;�`�K�o���0q�e��*#k�-w܀O~�ø��T-f������[���cؽ� K���_�ɉq��<��:|� e2�h�Z�S���&�����v9������2���YUje�&b���Kq�e�I���Wwb��Zp\��G����P�?��D�rIs�k�Y#(�a|d�h(�ϊ׳����\�a�V���p�{h65�|!(,�i��Cy��V�4�$U�Š �^Z<�x��w�u>������H�����Ͻ�Ǿ�^~i�i�$��굲L�.��\\~��(����jvu�����#E6���1 �S}��R�o8���ryE=�!�3�k��e3��@�bS��[��VuR���T�hV��������Y���M1I��f�e�Ӡb$)I�������5]hq�YRO�����yFA Ek��+��ԃ��g�j�E�'���@���R������SXi ّUHgF��+2���9,5k��H��	^�T�V,y*�x��3 ��Eܜ̒	y H�����x���f}���S?��;?�ǿ�3��(C���/��}�ڹ����Ӥr�m�ٚ��Cߝk���܉n�X���y���뺫p��Q���d�Čx��c%�n<�m���ٯ=�=3�����2�I�q(�S��c�j��o��:&�YiW���>#.L�_�d��a$?��}E�}ZY�F��(YfĻM��2���
*�%�c���KeU�[U�Ԫ�(/�P��vd|Cn@��'矍/lRZ*��\����`�@,��(���h�z��3��<;XLI�So�q��t���,��Ӏ�{�ֺl���8���/�#�Q��[A�5�0��?���c���|��؃riY��~(G(U����� I-��$5��VV��@z����V\��;��m㵙Chf���� ��D��$HN�1�L�󬇧�0��2����hCe �Q:	y�:p���ԒBs�5T��{��r>Z���Ã��^ga�5�q�1����B@�𣴟�A�,���5�Z�0_��mW+؉f�# ۲ ��B�����4o�Q�f��D����TDf?%S��@%�4������^ �r������%��U�N�B�'����r:���<,�Ȑ/�/}N��ړ��0T7B�i���Ԯ���QjR��d -<�5�ea�y�1C��`JN f�U��4}���Af���
:��uoTfb�E�t�ZH�ވ(h��`�i�(��RT�H[���z��){P���q��&C�ă8Ѭ�Lʿ��S�l�ƨD�W�5�h_��� Ga]*0�Z'a����C���}ݞ��D׌�s0�S9�>&Wl4k`�g�}-��PE�Vx���JV�b��s)�|���t��s8��	X��>���P����ҺjO��#�E�2ҰT%�*�1\%Jbw��:��D:��{�c�ӏ��ξ�
\w�ͨu:8|h�^��������\�Q<{����/�ͷ��F|���(�
	�_�{ �z'���o�����s����~N߼A��+�VM�t�pM�zbaǏ׿��9���&X_�~=n��Mz�t�޳g��0��)j�?~s�X�n�;�<я���ѣ�5^#�Q����2��ǉ��V��m��b_��t6m޼�s>�F
�s�>p�O�Zq��i�><3h"�WS���LNMa���Ԥ��3���wan��^,-9L��G��7q��oǧ~��X35&�J��������}O��K8t𸜿������F	�O[�_��w��[�E��6U    IDAT��L�V�H�rH0��f���^�KU��I�eOf� V8J�e��y��łƏ��?LR�4�
�s��qh���8���9tU1.�E�gS�>���n�Z��O�-���"�ϝ�H����I�Z=��.�*�G�W����7J�=*1,,�(�d`�^E4gm��f��S��u�Z�&�lD23�D��n:�x>���
b�rtU.��\Z�̡CA 64�7�.J��7!,³�B��	���:�y�S�g�}�M��_y�K'������S�!��������_��Nzb�����"A��ߏS����V�%P�vlJ)�NS�
'Y���W㎫��M�]���$FRT�hjsϏ�����K��4^�q���8VΡ�Z�J7i\0ʍ2��p�������e�ʁf&�Z��fMU������/���4�|F��r\v�K1�C<:f-�U�	�sQ0���@v����F���$�,Sqs�aT��X�0&���R�NJ�ȬSɀRY4�4��i���߾޷PȡQ�����
�ʫ�bQ	K�c�TBcv��YZ\�k۶����@m��E�1��{�.q�������N�>�̪M�D(Ys�O����[n�MoV��;�A1G���0 d�����CV�dL�Yvp�ˀn2u�8�����C}����Lф�g2�h�^L�=���`Y��u�<�sr����!�(���(�@h�� {��m΃�<��g0��/�+~��'WB��8T?
jHݞ+~b���L�gn���o���9�U$J�� ��LAA�!<�ISճ��4����fe��,lA{-��t@�Rnh��\�Nwwe�<Hl>�}��
NӧT��ЏQZI4������A?�0�0�>u�y�KT�@�a����JG��#�dR��g%�=r噅�P��/p��W����Rҿ�7)�h��,�C��@u�п%H5��Ȼ+x JΡ�ިJC�zL<!Wa0���{X�<�gә\ўK��BA��T�h*���Lz`bh��n��Y,��g��`���$Z=�k՘G��55��%�ϡ��]���B��Ẉ���Y�n�0&����n��1�����}N@��Ku:E���v�*����"�ڇ��y�n�]�z\{��(u�ؽ{/f�cn�4�/�_�#Ɋ4��4�c��7\q~��?�7^u	����2���G����G����o�[�z��ޟ�����ȋ�@��m��]XX�=�����Y>|XA��_�w��.l\�����#�<����,��@�0}�����,yfR=���r�|.l,^�n����P,..+���sߩW+J"���kar��k�ŭ7߂��ש�w���x��`���}�Y���˥,#υVO���W���8+!�Jm��
X�vJ{��Wv�k?��{����*�
D+���7�7��'�z5q)CM��_�����xjJ+ud���(��~�t7�r~����9g��e��� =���=9ڇĈ;,k.�������~#f�j�E.���Ϗ,�<��٬��M��p~�j�ш*K$��e1"ڕ:��2�k5�g��5Vl�Y,U˪n1�*ݶ;]��u4q�wT*W�J��`�?g�^�5(��g���s�����Mn@ft-:ǓÊ ��:m͟����f���_|�Z	ٴ)N1�#�#��	��zп�(��&�XB���&���릏���y�$0�����_}���W����8:~z��J_̀z@`<~f�J��7�j$,���])��vn��R\��8��H��T��IǸz7�.UyR1<������Ɖj��z�W;ʞ�3��!%��T\�g=V��G&��o�ۨ1⬛l�K��\���L��:��&�uX�a-
E�2&G�ef��L�'%�=5ɟ�r]Y��Q��Q �}3&�51��(.�S�e3�:f��C˃�\/���M�U��>#WՐ�v~.�:(���3M�6ҩ�&m*�C���2Yѓ��c�<���;w`f�.���Z
��L������*�l�:�0g��R-�}�64KIc������7߈����6��8����֠$�fn�y3��T\�(��E'1�?nCn�9ݲ���5@�kA�yW}�^�H<<��w�C�i�j:�ud�4��l��_��U��;0�<��k��u��!bWAN���E_b�8gP  ��J���C���Q�8N*'+h��E_�q��tMAJ2
���>�;Q ��
�=��8Y�ҁ� ܠR`��A�0*�载�c�He7>��Z�.r�N����$�����������F����������T��q��/��F]:P��!��]��J3��0 ����Av;PTLrZ���0�g.`x󪼅�`؃b|d�읪�*N��p��`Z�C�|��)�p��a�>)c�b��� ���������@A@O� y7kc2�ǭ�(�N�� �r�N���a��������6
��r����2��D�<���N�ճe%1��q'���2����a��s�oE�S�U�\��/{fV�L���q��?��|�z�f�϶�������������rӎ���w�],�T�w�~�3��{7x�;�<hj_�4.��L����t�������?�kټy���ࢋ.�SO?�/}�Kؽw���Y�\�����u��a��*
�Acw&���LI��Z���ܦ� ��L*e������:����pƖ-2�z��g�����jy_|1ι�\d�#jNN�����x���%�m�d{�$�_(�;�~
_y�;X�t��Qo���8�T��{����	#y�ڨ�;x�����*^ض[ƥRUH�i��iW�zUx�x��ލ�B����@��������L �n���_�%<}|/�\����Z_f��t�)�c� �Jۖ ��Н�x��n�j����+KR��ZmVZ���Ǳ�E��}ӇgQ_�l�By�ːݶ� �N���hdKV��rh�J*�E���- %p���Dt��1Lm8]t�J�#��>'T�ׯ]���?_�˯���C���`��؉̠K�;�X� ���;%T�pS�.��%��=��;������{^�	b��~��_}�-���_��F���0~:�1���X@ЍO�A��F���\<ifV���Jj )��8�&��sq��c�d��.
��8��,4�i ������>��s=�G7a�ƇM|\��#�F�]���u�ͬ���r�nD���:�8L.��a˗��:�Y�����X��u0Q6����e�&�uFÌz�WP�6U�'g�J�$�aMM�)k���6e��6V���������(�U5MMLh�Z���L�e���b-XF�t��J>���2C��N�/S���6: �Fž��c����ۿ�1Y�dL��Ǎ�Fn��{�~��3I3�����~4s�te�t��N���[oƭ�|�ʎvH��
%'C31�@R�@��#4���qP�2p�\P�-�4�3�T�(@��z|?PN,�f��APYz�̻te����=�y�)���� �d�ʸ钼b.��\���0 ������u�쵫 y���hU ��x�݁�߫!o4����t@��1v@��yRfT7\I#��?�(0>����v���g4�#�ۯϫH���:�!ȟs���ʯ/�J}��D�}�Q�&4����S�a ��(0P�8'Dz��K�N�S������7�ac�kr2U���M��B�!\OtD+�'�(���92��xuNk�A�@��di^��Y@1��G�*�&��e�5d�S%,��D���s4�����J��܇�D��y���M�����Eш�`,�d��ϑ�[ Y�y�9;$�Plߧd���0s�{�'P�z��"V��15���׶���>���W^�X1���Ә>t��%TfN Qj"٢�F[8ڍ*�e��ʋ�O}��|�~��������O��f�D��wގ_��wcl�<�����#>����XZ^m��O<��{�o��?�	\y�U��#�೟�,^پ+��5�j���?��n9n���ĥ'��}߰a�z�(O>:��$n��v�灟�کժ$=��G��7��NW_uν�\іFWM����L<���	�Y�J�lͧ��yf'��K�����4�1,,̡ߨ�]������IRڷ!Zѓ��ğ�ŗ��+��ɏK�V�"�c�C	S�
��O~��&�%�"-v�e�\�,�0^��r^p|Ȭ��V̄v[�ȕ��l��g�K������m�&�Zuʠ�M� 14���g�Cme�҂��v�$���%������m{��cOb�΃(��Dvl�U�왒.��g��h�!Ms�P�	G�����zp��>���Od�%ݻ0�����4� k��g�*��p�ƍ�2�����=J��8/4�Km�8��W4���R����T����Ҕ�O���ۯ��g>�3;�g�O��j@��/|����_��j'�9�j�(���^��^�l�챔�3�~������ll8W�s6Κ��Y��0��c�h
�\Z��&K���m`�t_��K���z�uh��$�:-��iЮ��0�|��L���6YPE���fO�C�Rs��߹�v���9V������2ҁ��" �9:V������R��0o�.���Ln��	<lr�c1��Rf(mS�P���byyI��f�9��U^^�ѣGU����f�ɚ�,�qm�;��S���>R�"6�s��0�RQ��l3sG�c׎�8qh?:���ǆM�AF�u� �����Pc9�e'	ތ���6И2нfɉQ\s���]�`!��ieJH��¡n8է"�˦3 ��:_9H,�(l��r����I�<�;�6����XB�CR�K��Zm�2��fU���?�A�Iy������V)Se󂊗�zB���G�P�C��ep�s�3IP����8�{@�����t�8m�k�E� v���e޼7@�$
�"����aC�1�5�Gʹ ������(EI���+
�e2(&↯�V1���O4C�A������B��&��ow�>5X:5p�Q���j�1��(���q��kX+[�4@�3��W�zj@��j�(�VU�����H��kũr�@%��8e��q`@`s�+�ޫcS#�L�����A`'*6�Cp�Lh�k5:7< �ߙ��9�<��l�!f��}���0���f�mmY`�ʳ���c� Fe����@M��p�y�KRD�����V�fѪ� ��a��8���Î�{U=�.���u�`��,i,٤�U��[n������+/F>C��£�{��7�=�����$�o܀�o�o���ذnV��ٗFi��cǎ)�$3�LJ&[�#X\���̌��;v�3��/��:�̳���_�2~����}&ɲ��4g[��<cyF���� �c�&Y��HqPae␉@j�s���"<R(���~7���2�����=�o|��׾�*\��K0�j�\^��Ջ��J!G`�N��jb�VA��D7��+;��G~�c�5 E���Q[:�{����D.M����N���g��M<��6��ZV:8?�.��8�x�����x�[n�!)�ʲ�TA)�1R,�ݭ�a��kC��������s��~�H�%=�� I�0���2�i,��JJB�j_}%9S���O�+䙡߫#�ĪH2��**�j���W���^܁t��$�0X�̤�S Z�F��KaJn�-�,2Y��K,d���"��i�q$ؐ�/������*�E��4/�	|O
6��W��L����g#�Jj���?�D1U�̿KL�^�~�'3�����>�[�ۮ������O5 ��_��m��Ͼ�߫�������Et�P�!�2 ��8�+�*E-[�/v�j
I$q֚���s��3N���ǑC#��X;��n"�F,�Cs����
����d� �U��vYv�/��� ��� ���уd3��i�F�)�q:�$bH�A30�1�W��!�[镁��5��R��Y�u繰:���k��o��r���D�Y	���H���P�::��s_�r�t�t$cciJ��_�W�13�߳R$f����N߂����<��΢��e~Dz�ˋK8�w?�Duz���k��C[�h��t �2C��@M��c����p4�Jŷ�N��x��A9$�
"��6���8<� $jhl��>_5������V��������FHPU��5��?��#i��.���U|�6�5Yʠ�������!��{�4�FA�'@����x�L�R���6nZ�oQv��sY��@�q
���A��5���Y?�ڽ�� (Z5��d0���K�Q�@�w��C��l�2d s��������W
N��H�p��-9}j�^��F�o4p����>5@8���!j�ʪ��#.���::_df�(��E�y?�E�	�i�)�a�f����������SA�n�}�g��e��2��������3�ȩ���3H�^�jw�<�ml#	�NV�@Pk�~����^���x���l�9�q���P��6�l��l6{�Ê%N�i�;� �ԜhuAUK�JUR">���o$&�d���6�ƥ�;��MbiyϽ�"���/���J���*��>R��f�H��@i�J#�$��v|����9�&n8���Wv����⩧_�=�4즛n�u�^���	�v�Ԩ�9�V73���14�5,/̣R)	̳y���4�;�|�=���>[�����������ܟ{�y{#~+'���)��s�&V.���l٢����Ǳ#3�t{z���~��~��{�������'�͇���٣���p�%a5��2��!�}�aO�,�f���[��M��m��`�+�Qa��0&@�����#�p㕯�o��b���{:�_�q_�ƣx~�~L�߂M�O7�g����,����߀���Ez��Ѩ��s�N�ܵ[~���}�}�/����D�A ߗ�f�F�\S�Ne������?L^��������Yk��i��D�K+JQ���hk֌�-��%�b�V	�^xa����aǮr�m1�O���W��=DK�cC�O_�$:!1L���/'TBZ�>���j�@�/Ic��9ؘL|H*�Щ����Y%E�>�{M��z*�Z�%H5�A8�ҴlIc�R���elX����o��c����v����5?Հ���������x��k�����-�p�xqvM��S��^t�we�F��FS�\v�x�-w଍�@��L���C����d�^{f���ן��?���$�����]�ͥ�Z<�m[��c���"� D�%�f_Bْ���Є��o@�2~��!�H); �0�c _.��;���3C�AzƸ��`��V"d9���.ҬC-��O�]sP��շ�Х�k����!���@@�2T�2E�t^�i쌳����s�����ѥ,�$�h�Z��w@��ʡ=��,H�Q��9[u%��+�
�"�H�Ǒn�$�7��w݁�'�u��.�j�sީ�{���c�C]+�Ԩ��+Þ
f"d�R7ڇ2�p빆��3�
�(7�  ��;�!
�¢��0MRM�����@�����4ό(xd@�>�< pz��U�+'N)jQ���6��s�nr���Q0����K̖m5�|n>���xM:=��(�M��Yց��7|��/�JD��6^��u�o�ωr�}O
���澃]+��~O��;h�&��(��o��`�5�c�:"��@��U�h0��g�i�T=-rW&:����`�1�r|?�fW]������Զ��zF��دك�`�5x��0�����O}>����ܪs�U"(��``�r�.��M��R1:�+`��f0H� �`?T'}.�\�3����{�|�_��<��~���  ��+���雯Y���g�7M�ȍ�ڦ�����i	�,p�y[�n�(N�ž}{D� (�Ek��kH�Sȧr3��Z�t    IDAT� �W�vr���{��<�͛֠Q[�<{��}������S��x�&�q�m����5����@i�a�RT2%������L2!v��4f�u��� �?�B�#����{��ź�p뭷J�����ضm�*�sn���q�
��ä���C(���7��Գp� }�Q��}� �Haw�}7��]8�s�4���g���������w7nZ���:��1t	4��1)�P���X =zz���v�s�B'WDfbR�k��,�O�������p��	5p�Zm<���x�k���
�cSX�q������+�X�=��.9z�;0UL!'� )@ֿ��3�<�/~�a<���ba\q�e�*󋀟ϙ��O��I.k=��{��߾�Y"ǒR���u���F�䛰ē�<�V�����j8���x�}w��ֳ.-�E����K���<�;��!�#�x"-�F�&cY]dRMUaJʃ)i�(���Ͷ�_���L
�d6�'e<�,165E�3�juT�a%3�U�|"ڣ'D?�$��3�>2�d�Z��:�]3ɪ>q��b�T�{��y�����b�����������?�dV�]�MFZT�P@@�8�G�H�bH�M;t�%el�"�,U���D��y6�{�}�`˨�&��&�9;HX����(�c�9]�C_}Om;&���Ȅ@�D.�3�F�_>�g��U���P?��<F�A�;P',�o ��ތ��{�TB�fǔ 0�Ճ�5'4f�c��.��	`�z|��\��('�2������N�XS�M,������� ���T1��A�Ar��1��͸���q��߈݇���)��l�f�1�� �oͣ�U��i6s|��7ʋ}ȸ�L2Aڇ^EP:P�1�:���T�bt�Z9_���<qL	�ȫ-A�;�3�����A�]Sh>#���L�� R����,��@M�Cv 2X�sH�zP0��ٚ�]�}��8�Ual����$y]!S�xs|4�6u�-dQ}����>�� U�@$B�1'�a��d-$�Dk�fzO��CE�(�q�س�|��=�qp����D�c�C*հ������q�P��"��r9�A3�Шˁ�_�v��<�*#���f����=(����Ų�C�S����� �:�'��̫a�8�X0�C��l�R��v~]���x����P�T��*��k�g{�'<�����R݆{�p^�ar��3>X�S�!��̽χ@�q�Qh����2�2�҇�������>��5����)(N�C�P�փj�N��q"PH����)z���(�\�9����>zᔀni���%���,�K}���Z���rh�*�B!C�_*G5Р�L������߆�gp�����Xc�ϼ���~[�D"�ӷl��o�7�|��b���۷++K��z�tZ�f�#9�����;3s���R��C����zTjU|��_����.�M�6�n��wީg�}�>��>���s�߇N��1�x�����O�Qk��nP��Aݭ���#��DPx��W����4Z����x��#�
I�@8�Mg���5���Q��$R�2��肜F;�Fi�Y�������}�gދ��Q]^Be7\r~��������(5[��_���=�^B'Y@:�S���Rr�{�E�v��/>�^�M �i!�ëx���?ܪ���uk%��*��,-
�z���F�$r�5�ù���������sa�@�b�#V��F'0�&�5�3Pe@������b�������y����\�blt�y�%|����g�َv�=�Eyh0@pO��{3��>AsGa�OA{��w��GTF� Y�CI6 �G'�Gn�&7nD'������5���Ń^�G��b��UM��k�*����=�k�	u��HJ�l�T��Z��������k����������Z!��?�ʻ���_�#�W�[�uNN��Rn���<zq��1��I$�%�֑��q��V��L?�D���#cxÅ��;���7�6u��@&c�G��N,�Z?��;��W���W����Bnb�ZW���i$�X�8�~�˘��,ОE<a����h02 ?�[w�@��3���X2���٬�P~�9 ��+Yv�XDS���#Enz�ܒ�c���5� �@f��>�N�Z@�_V�7#_��$�5�l�D$��T2�"��32���|&n���;�B�6}L:��zWҩ#�"f�ƞ�_@{��1�RU]8�e e�  ( ��x&ۮ��:J~���DM6��ȯ���܀7��V,�ۘY��l��?Z����+�^��$�7 Y���V��X� �@���h`ͫC?�( s�t*����!�j��s, P�},�d� ��B��%|�(4,�FmJ*2CB�fꐣ(�3�N4hg�������A��ݰ�ҞϏ�`B���*<�ςF��z<��`G��eC=H���{*�gN|z&I��H� ��v���O���p��P˟E�~���:\�3:tQP��G�<�9����ީ�= �A}'��>�B����D�B��d��5��|9�3��r��,�;Ѡ����cjOC#?�N��z��v���U3�D�<�(ষKt�G�D� �7'm�<�T��u}R�	}8�Ӈl^���S�����y��(��&L���Y3�)v	�g��7Wp�IR����oŀ�j���eu:z�C����i�
	��d�d��*�������s�����2���Ld�oT����8s}I�6ԗס1����ӋI�������2����|�C?�׽�l�����O��O��o��Kg���M7݄t.+jΎ�v�q�X�cRY�"Z�:F�yL�E����٣ؾ������>���{1�<��~���Cj<f� �D��G��׿�������ʆ?��������C�j��׽�BI�~经((au`|b��{/.��lݺ���K�teig�}>��K\��+1�Mb�3OcǓO"Ѩ#�
�X�y2cy$ٷ��{.)2�4'�JS�&�^��r/����S��ӻ�a���Ǚ��N�^w]s9>���cj$�t,��fS����l}~R�	ĲY�Z�u)��c-��|+>���ጩ�<Z;<x�������C�I�݄hT��F�����U_��J����TVA ��q:����)|�Fq�6>�j�� X����ZKKh4˸�����1\x�vf%Rx�����|�4�1d�􇠐��2��M%�e2'���Q݉XM��K��\��1����8�6��������g3X�k4{xz�)ٞB1�U@@�$bVU��+��� ���įg0A)}:=s�m��~"�����c��*��W��������ȯZ#6N��B,͛1��d7�d;����5��]�Ѩ.����N���#���+��{ގ�]�3�Iv��s.Ymm�1R9�����ކǞ;�fb��I�i���҈�g�����kO�@��d�"=r��Z�V:2��J����C��G�c�gSoD��E(�{m�J>޻�	����%(eH�P��>�t;�NV��I����Б�d@a�;�&���nh��� ������p���̎�.��o~;�S���14{��N�Yk#�Ob����
�l@j3jg�BG��F�(��}Eb58i�ׁ�������U�^�����+n���|�YgQ�,�vW`�,��}�T7 �Ҏ�6�5{,Ȱ��x��2�N* e��P.�S�V� ���#Vg�	��ß���U$(w�ʎ�T�O��D���cm���H�|�~iJʒv�5�7��f\j<��|�!�Mm<f� e 6O�]t}�9<>|xP=|���@l Lp����3`95X��d@�2��#���F�՝\�����:Z0O��]!�<8P\[h��VB���i4x�=G?o0�O1�6�?j�\�d���Y��Pɇ�K@ƿ�L�����ѨL�`lN�/E+7�����{�0��+K|=f(V��33�Qےc�Y��qp&�L��Lx�3��t�����q�̒�d1c�J*��ӽ�[����U���t:��O�
�w�^{-��������]#�Ҩ"�3H�̪~jj�>��zUЮ�4X8j'�25.�JVX@�	>O7:��)n��� ]A����[�;R'8^r��T�Uh-ZȀ���W��|�`�N�ҟG��P,Wq���\�z���u��)Ṣ���d�9��_U2����EN�.Q�U��\S��Z�޻��W1z�Gd!�WEl���}Uj��-����a�d�������	�t�|TJy��܀���	'�{ל�s���9�H��k�nt��#A$��T�l �N��%�h8  �(��?Ћ�;�������k�b<=.�G{===�D�׾�5,^�X�¯~�+����_�"�;�8��������_$��+V�����[���Ѓ�n݊Gz��vJ�d�����?a������FT�i���(9aVx�x�MR%�x��â��^2��p�qo�]�;�a����^�K����u�����.����`֤���+7�A �
O8��"�{�Tp�-Kq�mK��T+d����bՆH�3�`�<b����� �=W"��r�פ�ڥ�ւ��|���L&EU�!���"?���k�����l��@�r��	Dc!,^r)l�P�x�o޺|�q���*�������Kv����d �s� �hT�^��]���Lܫdo��H�xc��
��*���h�<��68=Ke��'ஹ�Y��6zZxi�V��А�Q��C���[j��y������NJ�k��V�娿����\����s�~��}�W����n��3/��+�����i��\)'%�/�2�Q�F!/0�4�u�ȍ����D�\x��Xv��8��)Bw:9�������ۋ��*i+�X} yW3�Q6���wU�����+@` Uh�R%�GF���V���SM@j�-I9�l/�&��d��c��v�QYm�UL��d\ܔ��r3��]Ӻ�: ��`�������A��,IP�4)�QPj4��!3�J�RY�k��
�5o�f/�9��@���:2���ɷ+Q,<x=�w�<6���=���P@��S��K��-�𡀠�I�M�T��8����8g�G1R)�o|�^r�`��κ��__���m���ޘ�Ӂ/��)`U���j��'P�CY�͋v:H%ʪpX�E� L�O]c�+U�(\(5(�3�))熋�Z|r-��R=J�}}I��W�%��AޤZ�n�|�Fŀ���N��+��t���fإ��5Vp�*Qz�KY�J������P���<�:x���d��b��|X�h+ A��E���{t0Ը6 ��{p��[�Ff�O�� :��k�)c|�M��'�@&�{�;1�n]��c/@��l��<4�k�wx��
��@_o]������i�_��J���� X���."=�d�mFc��?���'��_'��z�B˞ښ��c-9_+��xu�������ӨR��(J��5�H7^�5�����\v@ '��3�iY%:N�ǩqm �v5�կ���l�u}��n9������y�<$�U*�P>A�w��Ê'����]�������\��+�-�;R�aҧ�jW,�������.����8�ϟ!��|�5�7�'?�� �b����sp��c�W�unڴ[�o@��@�P�����p$���(�(16���^�4�qߧ����\�t>�g�}<���k ��o|Cz	,<� �����z*~�_`�Ν��cWJ���^��M��6�1"p��Ǯ��o���}N�H��L�6�����K.z�xzw��009A>��X&���Pe'�o�y�ۭ�G�~S�>[`ˁ^��Ѕ������ħ�#�A�Z���NÏ�~/BL`:�(V��[����=�������U��������.�Zb�3I�Y��?�4v���{7�i��T�������z=�I�ȿ�
���TH��d���ߺ����W�8�:�����p	��N,��r�t�M�:m� ���y�������|�U���R���%�g|}6���Y��Ĭ�QOȩ`E12h�V�(�!��j\����55���"�/�wL  ���O�F��U�Y��V	����"�XƤ\��ZH�3eP�jI�҅�0s	c����nX���|避؞�W���'ox��Q��)�U��Q,唙�u�~	:�.?���,�.��ƙ�,��o�����Ͼ��z��fܴ�:�y�	E����6f"D����@?���> �߁`�$x|�*��LTG���1е0��j
^3@t�k����Yge�1��h�i��q��R��8���	�l�l���t(�-�|���RK�D���
��Ck�.9�+e�d����b�%�*�j�%����"�d3�� Ȭ���{/jUf�0��'M��-��S�E��(��2�57<Uj�
�{п��p?PʢZai������}@ͷFFU�<�B`s��f�PY8nf��&�}٥bL6\�c_o�,`v��cQ�dY�2��iJ����jʑ��j-�a��4�lxSp�r+5�b(S�x8,Q�(��"b���]�|��;8͍BaQ�S6�{��E�M�C0���(Lѱ�(1F7MQȨ2��+Y��)��x�񘌍Ȳr<,�7�f���
f%��Z��J�˪ZsG^��1+��փ�������4��h�����B ��j�Q�xk�}퍀ٚ?�JX�9z�����U��D����������=�����q(5��9�Ϩ?���֞��_O�c�ԃ�z���~]-��'ip��Ms��[�Z8'8���l5��e�Ys����كi;�Ҵ<i@�9>�"V����6`��]�ܒ�U�~��9$�y��A+��ԥ��`X�[{@>�����?D']W��ϊ��%GZ�~��2&�S��� E��,�:���fz���ԥRQ����R>g'3fb�}��v!��'��i�$���?��
E��Ѓ���QB4���g?��fu�E�
8�z��: `r��s2���j\t�G�Eq��A᷏���μ2�T�C�nʚ�rH%ƑI'1�Ak<��}������eĘ���;<xPѿ�n|��O�ꫯ�[��!�a��?�y�~�i��~����ᮻ���)���/HǊ4����J���.|��JɀS1��	���q�E���`|�z��@��)��e�N���w�z������_��C(:C�NcKW/��;�!�����#���(�#g�����/��>Nd��f~��3�`c�Tl|�y�A|l��Rˮ�_��.�3�ٹ��>���%�񩠟 ����cLDi0�ְ�����/ �� g�%.�J��I�]Ȓ~�X�\yv�K���4*Il�Fc`tlC���5Eq�����n�/���_X��>:N�vQ)��U�7��䭗�¦)�A#�DJ��D�uR�]K¨vT�v�ܤ��u������� i?<�)s��Q3�(�0R��}2&��uIs��,��, Q2c��A�!�RY��Ҝ�-+n����|w�G��>���?�� A�Vs�����7V��g'y|�CQ�����Xn_�P\$/K���*:[��?��]��ډ�^�=���E^�s�>nO�	�jSE�7ǃ\�����6�5�@t�m�u��7\+�[H�k�k�۵0��d�vS�F����[<v+X��͍�j��MqCU�j0��Bu�ˡ#\�n�$�޿��ZN�܀ٻ,w��O����>,�e^*�=>�k&}�45^���X}��ұd�9�ep�PU�
U63��Pv"�6�^�ϸ =c)�$�֜����?��{Q� A� �, i���I�����{4�Ҋ;XEa�������«c��a�Cp[Mu,9K���"�@��	7$]W�؍C��oVah�N Ţ@0��~U5{K#�ڨ�Z�`M�(Z���a%�h�F� ��}�V9UKd�t9��P(�I�Df    IDAT�����z�Nd3���!�~�wO�� �5R�y�(�k�7�W:�E"�B�U�	ʫRM��V1kX���X��=8�gz�j��[�q�s�r����1�;���W|�H ���{@�N��uP��5���A�$�@U��s#���^{�� ��@�׫	{ n_�����?ĩX���'�����/���0�wZo���+-|U�8X���qB���fl+)R�UUm�	�|2�Vf����*�!���@�}��sU�_�q�ԁ�'�C�-j�l綀_z���P��*����x��ړ�E�.K.���]>'=a�>d(�&��#� �ڣ��5��@ɾ���\�CQ
u5�TF���h��*A�Z�@4�G��,��0�������2p�3}.="J4'̞��p�x����"
J&�F	꺻ੰ��D���γ�|��7]>}�-؟��٪6�{��6o�-�Y4ބ��='�r2::'I¤����I�����8.�!`��b>�B.���~�~|�_�m�nA&��O<����[��*���=��ƫ������{���`������?��N<E ��W����ҥK�5^ye�z�-�����M�$���?�1.8�\8k�ݍm���,a��$S�H����� )"f�N��"��/ol�%'�ŪM]�O�P�z����fQ�&�����ӿ�Z�!E�\���l�o|�v@ �5NRZ=H�F�p�W�s��/�8�s֬|�w�s�*��ʦ4�O��9�󌒡�՛f-�^�Y%�a�����)�����x<���ף̹�$IfQ�t���( ̴S��R-a��.��������;k�n��o�޾ax�ax=a��&�$J�ʭ�C�ٌT���|m&Ԍ2���E��JY�+��ǂ"[����O(��ˇb�	�/'�_�PLOG��(R�#��M4�(��L���h��y�,*m��/J��Q����ӘN͉���������+�]�7^ٷ���G޼��U�E:N<nfN�@G<��#G�f�&���C0ގ`s̪R_�|���h��pڱs���+����ޝ�E�w��yp{x�J�qp3��4sD�:0^p��]xm�TB�j� >��(Ù����qd�@qHz�Ϊ��۠��;����!�(M�ϭ,�ެE\h
00BR�R�ꐘPn�9�*	o�����i%��fXI��5�������O�TFu���C,��\d�6�*�#t�-W�(�0�"��+Nۦ��EK0���e��I�_�B��1����^���
=*��eH�ҢB|8 �@�?f�(C�6s�������A�� j��fa��Z�@��2հ�SYt�=X��x����Q�KƝz�4na���q)�9q���HT�g�^5�|�f�Q���9:��k�ӓ�X.#�ɠd$����)�*7BQ�`��ʬNΨ�����21�d����L���`t,�\� 1��73 ��'�,k�'˔���@'�����������u�&A��a�����gR��T��%��ց��\�k�_
,��2���	���; п�kک$�5[7�kd�u���uMg����RY6@Ŀ�4�~�r��P���������_g����@L�^��4�H:8�����o�@�xJ��
���\�ʺ�Z�F�%f
?����B�]7�|nT*��eF�� k�6�,t
H����jݙ2���S�M��phpD�#~�:�1�kTӃ���ާ�X����O���3K9A+���j씲����J�ݿ��fS�\��;�{��y6�UʤY�~.'{�hԙK!�sbfG3zvm�;/��R:���	�)�i�����V� ��f ��H�\ɦ{p��%H����^�f� 6�kio�9瞋�O;U�ž�~��Cɴd���cB��B>�Z��������� B~7���/��;nE�P@��?>(�|f�ٰJE!��Ħb��g>��s�Y��O�m[�J/�H�='0����q���Ϗ>���$DBQ���1Q���~�s�:S��=;v�������~�%ǐȤ���2�]vB!�97ʦ4��H/Gk�O���,}��8C�NGP,��2Xr�����,���L�xk=����iW�M�t�Da���иo��j�{��?���~ ���QI�Q��lio�`�
JvY�I�&	0H&SG�x�5%=/����Z���I��V%��%+��t�kX<Xݲ(�����SV�Y�Y��s�4$SY�B2����W*=J�z�+fQf�i"��6�������rtKvx���Au�LN������<�n7|��V���n?��fF���F�v���$�N��l��"�&�r�Y�
�8]�`�Y�I��@`%�+%T�bg���;�^���q�A�������*o���ɧ�}o���O�:e�ҫ.�9�����#��x��W��K�a$k"��	_�N���t��ᦏ]��O>A���n�X��υH$$��	����i�T��(^z��W�E��O�^�M��P��al{o9l~W��U3�Q��^�ֿ���dL,@�!J<�T�]p�C����`�����2C�HE%C��{��'�������$�l�ڈ�"���鑅��H,�q��ʬ52y�uZ�D�-�e^��U�N&\0��iL�r��s�iM�+��	w�g,Z��g���\	�C	Y1�v�U���ې:r ������O�)�����k?`��Ԇ&R�8���@���RC��ٸ��+p�%��pz�^�ʎi� �iK6��u��i� ��l�ͤq��"҂X�Q41f�yؕ�m]���u"���Sc@�I��r82�GWSf%x����"�OQzJ�7*������P��@�IFܡ�M[Ϋ9�U�J�T����8� @�	��	I�t##cU�bYmX�>0б4�	
���%Z7�����_C�@rBSl=Pѽ2��A�~}�l:(�5��ve|� K��`\*D��^Y|إV�"��NS+��E=X�SI{f]��6@�_S�7);���ؒ�����v�Q}p��������0����-�Dm�:;��]�� {Q�^ �F��Q�T�t2�}S��
�
x�I��9 {�~���[��AA}|m=/���ڡXUt�c��V�'�Ru�c��T��Y}V^�)IP��$`j�����؛�uŉAw}��rҶ�����7���+@ ���\˸[�
\'�[��&]!_,�k�����
���R9�������s��6D��صqV��U�@K[��f��,+e@�b>�a��� G16����8|�7c�����y97n؎��a��D�b�ٸ�+p'bd|Lh>�Cê����O�+��hXV��J�A:���� �c�s�(�=��3Bb�����Y�믿^�~��Ș}�K_��\( a��}���K����}� ��;＃-[�Icm&��ף��	'�����I'/g��[��Ï`����Lb\��Ц�f��O�4Ebf�墘��q4w�Ĕi��:�ؓ/��U��|g$*��ύ��_��v��J���������G�����ʣ�L)O#�֖ ��Z,Y|���`ӆ�8rp?��	�Vz��?�뢚�CZ��129�Ƿ�G�=�	IVx�-� ������r�հ���auB*%5�L�[�:>�R��|IL�(��~��Q�Q�	%�Ru��c�
��Y��ǃc������>�T���Wr�"�C��~&}�(���]1ӈD�h��.�d�be����H<Uf`ON���IB:��=�t^�,F�*=�T���fe��.6���誰�{h&Y�����m�_����rɡ�������翽�`��ϼ��u��|f����Z�g/섗m�`��#x���x��5�𶰑�}���_�#���S��ߝ>N�7c#9$F�Q!�M@���d��)�%"��mƋo��+�u��i�/��ׅ�p�t�-�c��+p`�{�����*c25�U�r+N+7V�|��v�ߑ)^w�e������o�f4�N(�����UF�jF4+2ai�!lf 5��jb�����L��+��L�>5��C@�� �ڞA��:$xh�,]~�x8I}p{"˚���p�Gc�	�b�TA�H�q��cGz�g�z����:�Q���/��L�9ĭ�hq�~>^�ਚ��sJ%�3�oX�c/8�G1�O�Iy��H2u6@ wͪ��hP��M��ۉB>�1N�ba��Q���ϋ&�4�QA����:puÔ� lim�8M����L+J�HX��,�$�A�BU`��h��l�"1�п�eNQ{����/�	|.��.:C��=����a<��Y
7U�3�l��:`T�dQ)�/��Fy�e��IO�ζ���ؿ�2��^C*�Q҇�����C���xu0�0�A���u��R�d�G+��}M�D�T��mu���C]�=��t[����?�y���~,����d?|�ﭯ��]�1���"�kBe^Z@Z��x�J7dn��^�p�5�y��Yb�C`4 ���r̭_UŬy��cC=o��n͟��C} ��n.�Y�w��w���Pn�j���-I�?�e─�k��P�!���%趚�� �~�4���bq�sR��b�I�QsX�U:A��b¡PR���r���U>�T�t�@�a�>��T�h���`צ�X����pҸ�aɘ���V /+�Lʹ�jʹ�����7.��_��s�
e�{�ͻ����ﾷZ�=�Y�P��d��Kf<�h��J�⪋n��~J��Q*d�}���тo~�����[�
��/��_�R����s?s�g����_��ג����{�t�� F�G0}�4�ٻWn�L��o�Q��h�@���;�m�����:?��O�p�B�6oX��<� vlۂh8�`$��i _*� 	��i�%�TvT���BЍpS+:&�@g�10�n<��r���:�er�����޻o§��Șe������g�޺]p�C2ߙ�b���]ÔIq�p��wL'܉m�ס��!�p������$1F0���<aҋ�#�y�*괽z,�y<�ċՁ���Jn�sK�N�1�C'�����v��B9G��ߏl�pxι�aQ�48�I]*�P)1{��q��8����IY������Y�Q�{���#�(�N����p�[Q���c7���/�k�?�r�t/�kR.���s���cf �ǻo������R#�"�I2I(�"=���T�#���L'�g�?}�͋��ͫ.8��9?>��
���G��?~}���?餓&}�֥8n�4��GJ���=C������]B-��QǸZF�WFGS �[#8���p�E�%BϐڨPE �c����P���A��E^<�����TB���uH��z����k��{��8��} ӯ�Ni�W%��,��Z�Q�����+����,lцt����X\up2�X��1�:_NX6�����a]l&�ld��\�L2�&Q<�j��4��c
��4�t#}EQx��"�E��a+�]�d ��uP�߇@�	Y�	_Kλ�*�Ι�d���q.�b��pa�o��|�ܡ����D�ʋ���?+A#0PJHbe�Z�?�@��y��0/�<{6���F�p�Y�=x�R�sK���&Hj�x��r�HM������(_+��
�
\�T�v�L���>tv�#�Ju �UyQ����O�����ٜ4R�Q*�����8F��DLwLVg����H&�+d�lnmJ�E�.(�l*��`PʋMC���� Z�!�7�X�����*/ Q����ټ��M�p�/�\�2���|e�@WQ��ݟ6�B��VO��u&��_F�̬����������ZʖA�q���� �*�%�81h�5J���j�r� ����:e�[��4`�r~s�Y���v0���b\(n�<dT��末D��۳=P�`V(� 3�{�Ħ��:3��ف�=p�vB�+��"����5�~�a�,�}ph5�r���F�7UD��}:�mץ �RR��zgl��-M閷�����P��	r�j26�*���%_k��=�A�
���ʒ6#�f/�Mq�I7\�L��w��2�5/���#U���h�Q=�u�w" ��%Vy�{<��u�=e����5,>���r��T�.c;�+Wv����3�a鱂Y@{S�7��lĚ��B!�<n��@R!��v�^6�^ǆ��p��W��eWa�V	�X9ٺe7��?��W����9s�aѢE8��p��A���!��	��X2��e��l�cE�	&�JH'�̩�����m�n`������glݾ]UYP����.�{v��K/�$Ypҁ��n���U��ob�ʕx�wd��OA$��0:<�U�Vᙧ�@��z�g�'?�	N:�$��|�������P7���e<H��2�pϘ:M�T.rF���D[:Q��1:X��o�ƁC}�DH�,#�M`ʤ|�s���[���m��pa<_��o����}�v+sS�M!�W賊��(.��"����o�6l۴���ړ�M�4V�MQL�2Y��6�2��h�ƵL@ �SK�G�ΐ��j�[�J(���b��E�X�*��$˔��H{�z���*�s�J"��{P��T,��Dt�dT���+���罠x}jd��L�7��5,��b�"4~�l"\��xg�&<��cش��
��5�ri�
c�����/��>'�\��=���Y�5��|�K� �ES؋�o���l2y<���b�F��J@��x�%�I)j��H#9����~�*j�Lv������oc��D����" �����-������={f�e矅k/�Ӣ^���\e�7m�����AlܸcT�-��!q#�ᄉc���������Y��1�0�����Ǡ��B�@���ӯ��K�m��k�?�*��s �
ý8�s=ƺw �>��WL�(r�<Y\'*���S&���T�|d���/:�	Dn���I	�F ��!?���E.9LQ�	�AO36	2�N-z6��#��	���h�A�2/|tC��&�����G���������Ç�#T "G�A&V@(��׃`�+�,G�H��xq4O��ؔiwLA��Gɬ��v�Q͗л��{� �{ ����@@�t9l:���kT�le���SYMa��1�cٔ)�J��L��Spŝ7��Aw�$i�}*�^�I�l�)<�Z���G������!&�0�py�k&���!����"�<u
�Ѩ�:�BI� _��R�P�dJ>B㠜�2+  Hԥ^��2��\R%b�����}��i�����rFYއ �j{s��C�M�(p��cQi����S��G%>7_�K�����>�"\�LT.a�@�@�G**8�B�E	�SΖ�:խ� X+0IK�=���FQ�ӲiVvH{R�]%+N�t��������dS'���
+ ew��)�T/J�Y�ESat����t6!�{��=��a�r��-�L��$�N�:3S�����u�1����| ��)�O����y�d�P���A������� �hjV�e|�A���s�LY�?Ng�c��ov�%����:�ASU&��y	֩OoZ�գd���
٠�	-����x*K���̲��c�iM��2��OUV��RU��c�� 5���DSo�s�@�+��d�**�Ȋ�{�
�)���4�s�a���h��� �G�r>��-4 � J��TG/�*5�O��i@���h�[�M�����T���~�̬��g��XUD[u[^ס��u�SVBK?>���O h	���b��Uز~��4�T���Gw]1y����uLz{���%G�Ĩ�wވ�^�Y3;P6iz	t�9�o����2�ך�`>ο�"�I�Sғ��g�x*��є4}R�M� ��YܫG�N�a��)��׾�믻J����xC*]���՗��gs.���� FGǥ�{��c�,��?R8    IDAT�d
��Gp��>I ����Ta*T�IIա��e��y���_�+wܱr�����~���A	�3�������mm�2��p�\Z�^sG'�&�B2]���7bժ-�+���;2:���Zq�7�s��>WY��C�4{j|�%t���A���`�, ��i�/Fq�֮Dz|D�P�$���,	�|6#�8h��0� �i�h�J+ܬ>ə/g�j\f�KW�<T�s*+=�8��t"-��b|�
�����˓j�
!�X�I�!Ǚd�"Y.x��*�kJ�`V\F�d��5��x]�I'���K.���^�����d2a�7���݇���/b�Ɲu��B>����� #@ܿK��?�1|A�{h/��6^[�c9� J�fjUMA��e��ꏜG���{ϯxEx���\0.ʗ�DR���c^��C�q�1�>7��3��2���|���>�_��ܾ���J��W�Ҷ���z��n��鎶����8�/�;̛�	#�G�d ��a�}��]��7lŶ��H�5x�A��B(�y�B~�}�	�����`�L	��팄|�9g�Y1��b8��M��ċ��Φ��6M�7�*�-l�:�{7�F���H�'��|6�r�D9� g�/A$߁D*�Zh!kM\f;t6(�ǂ�HX�`\x�Y6�
��?J���M�Ur�<homF8LC ����B��D*�#��K���A�+(kNx��ʀQ�`�������S����`�����l��e�O�7�D���^��5�c�bF��; ��1�̠���C�D%�q�C����� �\<�7���X��hu�s�<��_�J�I���Í�I��W�%�0�C��ȍ��U�Ŕ��A�	� 
yVR ���U,�H͔9@���0i��l���5��hT�.�,�@G�I����
E�ۨ`����Ȱ4�
@c����}<\yH0���t�=�0�wQ7�5��S]e�U"�9�l`��HY�AVJ8GZ��:��-͒�Q���Q�"���àU�r&<�vdK����oh��|n8�
璃@WU�$ش���Kc��-Ҍ�z&��8:*z(�[6D˚fh� f��M�0�̡�*��	5�O�>�&7� �@2A*h�3�" �T {�V�:�b���%;�T��h�V�v�&LD�6@��'J�U�
��<�̸ζs>�y��&ݖt�r��(~l�&{�(T���Fs��q&�8'��M����С��G�_�~��[�g�嵺�l 4�Wu!Z���_a�M"Г�](��K��WX�6�"�W���`g@ =>N��֐���r.�G�,��~Z*%s(FGl�'��`��E���G��@ $f��Z.�ټ2c0�c%��t��N�)n����э�Z*Hϖ�5�f�Жs��O�y���>얊�	h�9�[�(2}�X�����M#�sP5K*o,��^�ω��^����G���^��hP�t�����L��Z�׍��Fiz&��E�YC�߅�[�c��u($Bq������T��)���2EU)��ZEzlM!�g�І�Om�(����[���[wx��y��q�1�e��9�-�� �I����bT&��l�d?�����6�����ŗ�Bѳ�?��_|c��r�/��Ĺ�Ԙ�BU���7��*s�!

�<16�b6�ϏX�>����grg���c�ꚫ0k�ll۶���a={�A���{JR��`9bʤQ��Z�v�x3��Y�@�o���>��\Q A�QC��Cs$�O|�&|峷��)�{ ��CO��|��FU��k�J�ժ���8�Dg׎-B���#?��ah�&�sR�L4�JonRB&^U�֪WL���d�%�H���R{���(煇I&H&�]Nr)IeE�����@���^�}E�n7L�zz�HU$�y�၃��e�M��f儙Ϣ���������߰��"[�b݆-X�v���H�
Ҕ�$A.�@����k�����O%��f��}x��7����0�Ax|MR���;�ُ�o�7/:բ��V��'_zc����6w�� 92"qלAIx�r�ʥ�k��@�D13�_0���;���;�Xz��N��=������]��s�����ⶥW��y�н6mێ�6�z��h�x�+�����k��s/bϑÈNj�ɯ���%Kp�i���)W�D,PZ�LDs�xQr��Փ�CϬņ=ÈN] w�YJ<:;\H��o�6TJ	̝Վ��?F��=G��uHʌ�XӦMA{{����z180,��֖v�����U�RGGN8q>�%�ɗ������=`��Nʓ��/����Tu.�f���-tV�RyZ�S�V�u�
�"kGQ���L�ç��8Q���g�w�\�_d.+
�x�U_�C�bf#
���Ș�dS�?��7<���Ad��s2;�Gs�A�#���g�6���i�CP�|( ���
��m֔��|JXV�u��-�pf��_�@hRθ�b\r�Ȗr��h�mwW���Яh�]u�Y��k�#@��`�R-	��ZGK�ڛ��-B$�Rp&W���|�9<(U*��@>�� �ĝ�� <�@��2��8f�ع���M�����l�w��b�TJ���A9 ����V�^UWl��V �9���Y*
�i����$������)�V�` �M���s��7B �MH����GG�L�EQ���( ��@����H�_]*W�Ge�"jR)�&���T���(eR8v�\̝9>���y������s�A�^��M���Q!)�K*�B���:��j޶g.e��������!Ki����Q���с���3h �Fϑ!�z����������U�;B����I���/��9�`ZsK=�1��R%�5���Ё~��c�Y��h��r�x��6��upi��`?'�VYq��ȰA���2xƩ�aHRE�)ܒ=�������g�ܩ������2��I��G���h8�p���U	u�_�����{R�����qH��Ũ�_��P-���U�dg1L�*?�
2�ŵ���(�|I}֪���a��*	��A>�JB(�.V���^����c�e���cI���������ڿׁ�}=�^�S�)�т������+ȭ�|�Y��UA��ܸ��mB��G�RQ��)��Y��\N��>x����YC:1�X��O�{��r&O���H�)����?b���ȗJ�T|�e8��D��k�.tuu�Jl�t�z{�eO���j�lp�`<1,����׾�E\z�Eb<��_�۶퐽�|}q����J�󜷸쬈*�,�����228$��'���C�&FG�Q�����ԩ�q�u���%�1::�z/��\^���E�(9^�`D�\.� m(��1�N�ǝz&Zۧṧ_���(̊Mmm�SծT@<��=w݌��w'���3�L�Ǘ������Ҥ픀�r�wV��ڄ�J�P�^��]5$�b�%U�{L�X�l�N�v-�����Y�0�6��B:Q>]�}��)�E㴢���^��!�HL��:ax*9�֦8T���9��+�e�9X�0�1���1�) ���0�� ��I�
"� ���;��1/~��o���?���0�<���8xh7I��}{�l��^�p�b����� �S��������/aWW?��XK�a��8��*ܾ�BT�V���,#�
z�Sp�È4����e?#�Ҁ�����>��5T�<������-O�v��������~�@�_^~�;k7|���t��`.�Yv#N�?�֮��>-h�K��.D{P1N��X�n=Vnڊ-{�c[ݗ�D��f�,��%X0}
��,�!?*EEGa�U� <��y���Uشo�����!���qM7�����&?,���s���ְy���׋H�E�,��0�шL��	�(�G�/1����|.#�Ķ�	�X���o�;�~����0C��**I�0|��8��X�����'�[��y�jE�јEc&�	&\x�%/d�L�������f�l�I7G^/�3o�Xp�OJI�����\�}^W �p�`X�p3%Yf�ܼ��7�� |l(����{0�{��0@�Q+؞X!�� ��:�WŪ��Nv�Hy����W�D��'_z�Tr��\X�!`ҁ��QVL�f	����P���L]�!j
�XΚ>3:ڥI�%���C=6yU04<���Q�,�pL��l���k����	U��Ě�̱J���J9@e�j�LOdL�JTV�(	(��dd,�< �$����sf;�
�3A):�Z1s�T�#aQ8��3g]�4���������T�"���Ho?zz��&h�Qq˫lӅE�#��R�� 5��
x��dl*��id�%G�������!t1�,��pρ�\���#�;_(*
؊��/�2�/��ɸY��:���k�q��	 �/�jR�L�jq�R%I(��)z�|�V�Ipf��
��z�ϪQ]e{EfN���s�L�dS��Twx�%�縋���~yH:+j?Pcbʚ�w�ĥ�g�4#�':��A�4���@I�@pV	E�cfV<]H#b���!�s�O5����'N�4w"�H���MSb��ժHp ��h�3� �R�j�[�4��ɓd���S F��|��4o@�H����jU]9�\�"��yU��,\{U�w|�rGz��X�._%Ry@[$�~�����l=��١ֵ�׊e�%������:]�2k�Y�lpBe�� ��:����go^��i�bd���a�Q�)���ǉimM9+x����k�z�{���
FU:GůGK�z&Ŏ��
�M%����Vܾ�JLj�k-�Ux��5���	��t#�70u�t,��b\{��Rڷw?���Fbd\�����'p�p�q�Џ�I���0�RsgM�7��5|l�b<��c�?p��[�k5ŭs�\7��l2Y��GV��d��6%��9���R6�G�4M&��r.2�L��ٳg�䓎�g�.�C���_{o��򹢼?�������� �bq�SH�Yxʩ�x"x���x\�XK+2���/ѐ�����L���+��C�bϞ>�L\�p�2�r�����$�xt�_\�k<ê��t��KPLO�m(�Erlx��|jr�k��U��``xhɱ�|~��T����I4EG[�P#y~3��4�c�è�I><����@*�5��Ba ��x#�d���Qz.U/��@q�Ma7��|�]��l
/��{�E�I�H�&�O�A[fSèXz�"���	p�Q���#��d�ު�x���S�2z��0sJ>y�Rܺ�"��«o��"S���HZd�]���(Վ� ��07<�(#�@�U1���p~Zg��;�_�?\vEO�\�˾���<��`���^����|��t�/�1��v+�8~.6m܄��ߢxg�s>�,Y����C,�_���C})���<�Գ���-���#�y�5X8w:�霔��V	^��>/����<�v!�1�7��LJ��!)Mze���`ΜɈ7��ylڲ#E,\x�l\�0��xXp���Bd���E�pѥ�	X(��G}زl��ln�67N4�����Z�c��n��-��p�P�-_ï��IGI��#����/��*&�QH����T��L˹�����,�H���
t�5	�yˠ>��(t��Ȧ$:�9D_e!=F�
R�#�� ��>T�Cҋ�` � �g�P�2d�Q�����/ p�T������s�"�u�E˲)6!�i��ȟE�C2�U��2��"��(�q�bzg&w4!B�B&-MI����!�A��U���p��_2��`�Q|Gr5�q��ԼH���
O<�8W����^�p�l�۫6?>_���ҙ�
0���Z#�K��)���K�K���R0�&VJ�y��Jp�JJ6�D$L��rK���R�`7��
��� ��J�is��Rf֜Ҩ%@���Ѻ�gX���4iG�Q-��q�98㤅�����B���̙�:؇M��Io���'V�fR-μP�t������:��gHu��ϩ]�>;�BT��>�9&r�	��"�;f�����˫,(ב
j-��h�3���-�xMǐ�p��Z��j VA��YT��R�:.S�G5�k�Ή�H�`#�9�T������5E0��M�); Pn2��]g��it��gd�s�0sJ;:�Z��ڄ�x��?&P�KB�=f\1`�@�,}��J�ť�#[(H�� L�6��Ύ6�����0)��@"�C"�C�H��$9
Eu?T�s�̸�HfϚ�yӧ ̽�,J?�({P<.$	�"�Z���+���{M�3���2d�
�� �,-�
ع�z���_+.i@�糞����>W5�G�/=�������#I�����E2G�>o#jc�D	�qׯ]0����h�E�`�dj&^y�Ily�=ᤇ�*;.���g.V�B4J0ƾ�\	��(�A�Tn��*�����g՚u�l�u@=�;'�y�p�g��)���Q �upP�ٯ�}HX�e�-�&�BZ������>�%�_��_<� z����^~n:���D��&�䇵�V(]��9V.	L��D"�L��S��7�GKKN=�DLg�&5!҆���#g�І|�6DV@�I�XX��fϞ��'�i�f�opO>�^|�UdrExA9S�VB>7>��[����+F��蓯�?��{��L�9�����*')�~Ҫه���@�f�y�g0�SC��Yp�yĹ+��:ø�]��>�c\�t1��>�������<�~���f����>�LS %��x��@4~SU�� �q6�N�N�3E�Je&�h��q�^#J�g���A[g���o��k����K/����_���,rE�_V%6s�L�� ����k/ǯ~�O��0��?��E�H�����Wb�� ��a��N�w筸��O=��<�

� 2e��D*"��֫Sh�NwU�L�I�e�Z١�ܔ��3�a���M����羸n����nw���ܵ�&�w�|lٴ���o�ko���g�y&�:�t?.��x���lH�
X�n#V�]���a�O���ŋ1w���
�����;dfn�n�xz�N��5g|*
�`$����Y����{C��
�{�4L�9#�$�n�B2YƩ��%�.��H#��@P酊܈�0��%�T����j�%}QaRV�~���C�&0Ţ����"k�[~�"y���S��Y?�Tr�� �<�Z˶����C�
7n�tƭ�J�f�Hg�0���j��Dx�S���Q,����]��~	�8�I��%�Z!���%��,K����h��z�@�6~UM)�HO��*k*���i@@!-��oE�ڳB@���B�"w���b�93�w�^��/<=��1�J���>(�lf6�7)EJ�&��˼U�6����ތ�������������d���b4�s6n ��ll*��R�,N�:�ESf�3�C�t���d9��Ё�q�~�1<�u����=c�a�u{<+;Z&}ǥL)�3P5U�@��J
�Ae!��,'ηP0����������}н�ZA6�G�d`,���h�DE��9�r�E���X���FD� �|��9T�)�]8n�4\xƉh	{ġ��w�-�#9��b��J o:�B�I�ZK[���u�u�!��ah�%�������M�} h�9�k* ��;lj���<]ACϚ�E���
�l��� ˣ��[ �`p��@�|\E�Q�/@��D-_L�@��(K㹮赠�G��h� 
R����YU�T*5*�j ���?�	|�
Dk�̯2��w�����Pɉ��i'�Ǽ���' b�/q���x�^/{~�B��� O���bQ-�Of\I�b�2+�����i)<TK��{�74��D�-�=�C2�.��q�8v�T����������)��I�r{ѵ��mގ��$�� <~�q�-����Q�C*P�+�i�X�ש��������O%y'����v@,�DK�@?F?G*Τ�J gɂZ�|�ƽV�9��j��$F*I��Ô��5�x�׭b�A�<�(��'�� �]�>������گ"    IDAT�G{K���2,[v%ZZ"���Z�v~����}�}������M�&Q�����T*�l�flH%2˪"G�䟣Vƥ��SO9	���êU+�u�r�$b`J�)gK����A�n���NU�cr��M.�}}����
�Զ�dM7_���H�J24�֩7��RFkk+�3���Ǵ3��q����ؾm�$���&�'+� �}w�����1<��
<��gp�w\xd�p(��9�JpddhH*�D������&̙5>�;�m�>/�E�`��P�N&�X1)[�&e|���G�1�L����E��RI<�^Rn��F8H��Z�L��	7��@.�D*���1��D�&���؅ޑ�&`P.����j�J��zǤ���#72�i�:�o|K��T���g��#O<�#}8ܤ��~��\�$n�a	����"_H�o�n���S �#����g�����{�3gM��?q��}�e���_�o��r� LwH�A�]�G�LV� ��4�)t@�F0S1���Mo�p۵��S���{Z��s�c�������xG,�;n��>[�t�x �wlCk�$��̚�������1ӧ�=�b�������9ԍ#���6�'OE����.T�q���J �Å���k��a� j�N�kn$Kx~DB!il�E�R������ǡ#�ضu7����@&3';UDڊ4�i%Eቒ��I6��`6$�-{=��g��Z��)j.6�����br;�Ò�'݈Y�!"F}�'�oa���1k��K����tbf�T�&��WndS����8MV.
RN��fP���:�J#4%�Z�j`tԀ&Ϗ�#u��b����2F�/{��l�.אG���H����àS1ui& �Vv��]��T�� ��Y4]! ���7]��?G{�B�����t	�+x��#@�'��PE$p��9�)�[����(����>�	t���t"�fi9�����2�adՀo	2�xhaZR)��(���,w(WP��<9�yr0���EM�A�
,=s�`Hh:�����5��5��\��eeKIߊPI��p���c!D54�C�%{P�eC��ՉD����dF3E���x�x��d�T���[9.�VG��8j�$�O��E矁���E���d��P�y~����Z}�Y�f08���T|O+*MX}���u]�
t5MHg��R�{A�l���r,J]4uE@�*0�@�G;)?��ld�2�:��*�4�IӨv�m���w�A� �j:���ܱ٘Mw|S�)]�ݠ����/Ҡ��|��̼W��+Ry�YM�"�jֳ�eU���$#Q^b�@jc7���0�s���لsN9���DɃ���ZIhM�B�*��"���(���
Z�Έ!���z��J�{2�L��|�Hq{�'е�G�FD�}�L�ufϘ��N���-��悋"g%��Q9�UY~>u��!7X���k6as�A$�8�Q�%����z�N��8�J����A�� �>5�Kg������h�״ =��\��!z��1�b��GQ:�uso�&i|.e����ă�ۥ�C!���U1�UMl\�>���"����D�ң�z���֖	���?2ЇΎ8��f�r��hmJe�������O~���!D�;
F�3�(���˜3|Mm�D�nV��p��=REktj.�X*�����5�d���_�ʒ.q.
����Ī/Ar&��,��=�t�� �.+��Y%3��aYdk���ğ�y�|�wM��!/$8�1�]��jFL�x��"_��402�m�wa�.����r.�b���޻o�W�Sz������X.������s	H���,�7ED��`�>���s/{�����,U9�U]����n�o	-��a�����Ѝ�����+�3f̔
_� ����	%���2�F>��x�N|�S�JZ-���ρa
�Vڝ^��ֱg�_����r-RF�@�����/s�eYy��>'�X9vW�[MNJX�B���Ì5c�,-{<W�������m��e � %�D4Bdh:wWN�N����<���%���K�?Tk�j��:g���������i4��i���:ʮɛ⏾�{��C���<���y���p��p�}Bg��U�!Ы������b�N��B���-�2�S����w��{x�����$>x�T|Ƿ����ͻ�k�5!h�<R0��'�yX2Ă��!^��k��k^��'����/�ÿ���~y8�=xr�o���?;:��D"9�p�G~W^�o��?����_BrdD!�Hid��q��x��12�~��X̬!�/!�7�h �N���P"_M�sk�Ï2��(*=7����*m����U�$��	�M>~+�iFї�? �!o2<t��"�ѐ4�Irb��/�^ (l*�۔�j��"I�{=��J�,6��/Gv-�S'�#��B.�VW��#n"���ك��A]o(�P$�T��@��E�Næ*ȖZ�$�;�4gBl�D$^;O�<u��u���tx�l�X�/䰃�Ӕ�� MK��=t���*���@a~hV�d�D=��ڐ��ҟ���l����9����@�]D'Fq���ù��j�
�;�o��ӡCw@z=42�	<زi�c�
,� n�d%�`�@O%�vׁl����euR�H����g���r�����P�ǌ�z
b~�1\b'S�gK��p�ף�c�m:���Zz9v/�-v��Pz�4��ՉV"K���JZ�0.ȼVI�����up���$�S��]����&Ć�bQP�R�|_Pf)�����h;|���̌����$?s�rsv��p��p��طm�^y�����-�Ud2�㎪�iP�B��]��S�ȕ�px86�C��σ�8S��y�,�&dژ{[��$�fraag�3�3�����=x�|�	[��3\��B(i]N��t{�>Ν�-��i״���.x-̛ރ�OA6�Jd���-r���*��!���[_O�y ���		?�}����[�G�c&6G�N�I�9�;�ض�� ��<Lg��\]�]==l��E瞅��0�lp�Ȭ��c�������溒b�H�g&26���H������>�GD�%-=A)�5��e+x��i��^����|�LN��9�v���&1u"t��¤]�D�K�^�ˤ����
y��^z�V�d�F���S��Aȟ�0�
ef��3��ƀ-�>�ٲ�}��0g��.7� ��?�$����~~���9��A�~�/�ؙ���A1
=s�K�G���HO�Y�^1v������T���a�	:?��%�>�d�Z�bq����^]��P�}�#��ǯ��H��U�<������L�,��e�٧�=�${��M#H��8AF/Hb�}�+�߃J��	�G�RB��F��|&i��2g3�V�.�Nce��s�Y���J�9���N�n�h���8%��X�~������<{�Ss�_������%j�� �ϛ	���zU�ձ��"����ib�܁�KU�>s�-����� C\�K�i|��G��;Bz��{�؈ 4�\��ଳv`n�4y.���	��E��Ԛ�,p��kbA�u�i)�\�z6֔4�NEx�{���^�{J셢�4s#W�4�v��XZ�G:��_�'\|���x���*p�1�ς<+w��l_����ڷ��Z�|�*M���T�ԁg�K�C�V1���O�����M�H�C?|�>�C,, wP�[��u:U��5|�#����Hg��������~c�q�����`?�3e|�oᙗ�C0���?�!|�}�"������ _���kN��<O��cJ�B��ĉ�'�'V�J��ժ�U�����߿�����_}��� x��顿��]��C�?���L�����} �]�Ǐ/�|�+x��P��x4�ljY��{�l�G�~?���r�DCN���BjE�{��p����h�����pa)ς��~�z�!����k�k�����p�� V�y,.���\�!0pR��~v6��#iT�*^8%ɉ� hkT���$٘M���ϡ]�� �P���B%�A����U�bi~�l^H��ba��m*p��A�`Ӗ����1��Q��E����**��z-;�#̅��Ö������Bj,��뫃e8"�::"fRzKp7/c��z���ώe�!S�x ���7�Day�ZI�v����2��k�Iov��vVG]�-����Uq���
�"e�Z��#� ��8�+qޕ�"[) [�[�W^��g�pڵj]�^��	l��pB�H��ˉd<��H��n?2�=��t�PX��u��Iu�Y 8tp��&o8�h��0����kD�4	O�YS�Оp�Ç	���������#$I*4gbgX�.[��(��@�
��3�Tʘ��C|c�@�Ϊ�N��J���2�� �brj�$q��)���d�U,7���b~��;��L���3S���̉5%������ٵ��>���0|h��h�����"�R���	V��]��j+�
��Z�֤3&'`=��y׍�4��L˔hX�LM)�d�LL��݆Y��	�*Hmؖd-��-I�v�%�UBH�d���mqL�ɭd��da��y<�h1Av�8���m̵��F´�SVW��S�KSr�"��x+q��ۿ�b��ې�����$^pҏ,�����X�����j�eMAl��o6ǈ�Nh���D��D��ÎM8��pK:�#2%DJ����3!���*%�J�~��!����,�DRe�҃L�(����p�I��_�S3�8rds+�Z�J�����8g� F�{D���Nq�@ilWa�o�^d���o�᥷�c��A���h�D�
$��p�z�p�Kj
�R���e\-?	��,ޏ�зwj��{�������01����6�݂}Nk�����]$0��{I9ɜU�Zwxa�t�o����c���x�����sϡV,��gM>� i�S2u�]NĢ%Ҕ����>��?y�JHY�'�|����
o�}J�P�zoP�B^7��_�abc���j�<�4�����Z9�v%�6	�jN8�����L
\0�X��<p��)F��:��gC�8�c�Гi��-8�5���`O���%l�gby�Q���gǜ�$�/đ[f��En nO���@4�X�� C�y�-����W,m�YX]��<����8�h���n~�gϣ�[����`~nO?�GgR�cA`�m?:⹆BgxF,^x�RA9�4)���yR�4�~�i��=1�;v��p2�fM�X�.��B��zC{��vbuy	�\��u'�굢��ս��@(�;��L_���y�C�[Ρ������l9_�QU,%���Y��� ��}7|����� �Ɲ�aa)�?*~����.R������ߺ����K�#O�P&u��W]s.��2�0�?�{�?VV��n�MW\�Ë�~�$����x��i�D��ϒ{��"z�t\^�u���('��n�b�21z�k/���}��<��_8=�߾s�_�yb�W{.Ox(���I\|�.���a|��;0���p�O�"2�(�h�0����ql��瞍�.9M'%��Z˨x�&/�t�/�<�����౧V���_EÝ@d`M��e��&����|h�+R�`'��W�<�L��f�j�Lg&��s^Ȥ�>�P��*e�t�j��*V�x��@�C&A��
fO���l�xx]/�A�p'Ǝ�`تc�x�K�!�7C�o�#شe�d�.��At�n�,汔ZC�
� �#Z�����Tpb�m@J��Qv>�H�	��7���Ǯ
9�Y�=����6������h��ͪ��88�h[����0N�2XxX�R5I��Y�7:N��LA�
�u�b�a��"8>�׾��})��,�4���	&���0.�$V�%+	�ߛ苅ߢ�*���a �l�4�ɕ�(D�%@{n�F݆$ȸHgʺ���l����7.���V0hm L���d�g�l\k�w�s`�Z��;|6L4����gI#;u���&;�:m8����k��;�F�x�ֵ�y�f�B%ݨ�Nx��ؐ84�t;�Ƒ��B���r:�t��t��1�"�u,�q��i��i�Ь��f��َ����~�=�0)lIC�X(H��K�6V38:���l	�BM��&!>����䎞T�����P;�5S�3Z�Vyg���7�p0�v�08v�ׂ�P�|�Z��r�+k&x��ҟ��yLWP*e���0�]��	1d�/���fvA �}��F����?c��F�R	�E8�{n����mw����8Xo�7.�y�R��u����<˚��i�2��Wm��k�q��ٻ&���-��o�	 #�` Q�PZ�햁wt��~��J�:���e>3�Z���o:�'OM	8=At]n�/q��N��G�TU�Iu������;5���}/�!��ŧ�<5��Y�K�C�u�7�.�_?��
Z4���k�Ju��99�#d�Rb6ɫ��%|s��?��LA`?�w�gְI�b�^��>�����ޯvqH�q�l�#�1�qR!
Z���޲бU��: �ĉ�ߋm��@��g���"�xnZ��d�<7��'�[��ݠ�L���[���?��n|/"a�|��ƳϾ�����ĉ�rq�:�q�a�[{}�Iҥ_)�9��(�Ѧ���X��f��H�Ϡ�&��>U](�'_��pN����&>)�5YD.D�W?�5E��2c9��4�,U�yk�l�A�ꬓ��=͸OYp��*l,�A�CDe�<!M��yv�M���H*n�X�iB��߾���?�����S�����?��9{�ܛ5`�����S�%��
��0/��$�ڮ��_������к( ���Q!�^�:ŧ#���_���"FFF044b�7>�r�%��ʆc��Ć$c_f-���n����o�&&&FP�t<#�U*Մ�hv8x�8�y�x�Q�/��.�ڒ�!�<s�\$�g��4:�/���q�u�A���܏;�u/�VJG��Dj�"r��
z�on�4��������O?�?�f�Sߌ[n�$�;�k��x�Q,,������]���㟽�{Ͻr�Z�P���1�/�|�)(t`x�r�(�ΗvL�?��.�q�M�v\�E��S��CC_���<���8\�`��ƍ�]��/� G�Ʒ����ȈL���$Kk�hS~�O�'v�ރ��?O��R!���l���ق�g:�r[��w{���x��+x�g�Qw&�@&H~C�dG ����l!�7� �hL��T#��

��xR��xr:3�q\X�T	�Df	�;hԊH��P/籶��J1�f�"+i�g����O���`����U�-��)-_3�m[Zӄ�h�́'�G}Ɩ���"C����ض�l�oى\���4f�WP%��f&r���w)�H�Ŀ��A�/u���a��MW�0��+�=nL4K�@�����N:�Vf	�S����*�d`F��c�9�&*a%`|~�9�}�Q��E酼H�b�%41��{�
�T>�T����g���>l���c�F���!�eV�З�iĤ��
�rzfG���H.10(��O�Y�䪺��Oԁ�r)�!�F� ��K5�[&�-�P�@/�F]�������;�C��*��@0h��� �������M7���D�Ru0�=�E#z�B����%�d���F+���HHd�Xȇ-婒�r!�/`�P9���j�H�Uu,��钿�,��Ψ��]Ă^�߽��َ���r�6�)�>7����x(��tczq��W��v�����.�Pm����5�%A!l쵓�d�ڴ��vw�.�dx#��H;Q�����Y��Q���m�s6�Cr�L��-M�䙰ҵ��n\w����^k���I��!���<�τ�k�����"y!��n���H]~~u�:̙��\���;�����B���p
,���򕁨(�� q)qbRƉ���U�̾�    IDAT����..9w��=���)���	~@�)�
*g��ȱ�Ν q^�}�2>�y�)�\vى7ŵ=�3���.��y0��cf>������BJ�?B"��[�ؿ{�}aM��$[�o��X�	&T�"������Lϼ�6ϤQ���J�*���-ʞ�zq���G C�ؾ�v#�N�m�����i������Wٯ�� ���b�1Ʋ�KC���"��ÔjmY~��Uw��m�G
NZ��6��6< ��:�6�vb�`?���}�Q�8tA�W]]q<��,���E7�.��V��l�>���w��믻� l#�;sz�<�J��j��r�n�?���=gM�%���y�1��F> %3%� &@ٿ�yEU�����j�
傰�:5�M1H/�F�#��B�((�'��������2/G�z�;u5�(�۪��RLn�4�����7�qϕ��h1��^��Orp/�H�Ӵ��`C�����4��ND��6�O�3�~
���C"���^ZƗ�~z�	�.���D�mx����`�WV�q��!���l�:�H�`�k�]@"G02�^��8�eH�l��l� �.�?�������'t�C\��!>c)5$���ra~V<������>��<�˭!�+"����GÝ�y'�����Po3V�D�Eu?����E$X�Z���@��Ͽ��o���<�G�{������p{�t�P̢V�` ������/܊R��ǟy?y����q��=|���-��QD#N�}+3J�a���]A<�ӟᡟ<��`1W�+< o *R8��fA�f�A^M��:t��\�����6z�'n��?}�#����� ��o|�^;>�����P"���m[��^��x ���P �y���@"�g�zG�~��QRJ<2`�c�G#��uW㼳v�C3'���Zp<:n/�nB�z���gq�xm� *]rt��008��4�"J�JV��pD���d++)Ʉ�{!���x�>-T��� GK�r�j�Z��%T�)8:e8�uuz=N���p�X-���hx�!���8���F>��ԤȒ1��a	�ȍ
���Ф-YrL��~��0�}7������=H�"],ci-�B��eYizeA��d��(�,!4�pJ�P�	�C��Ȑ�H�ɗ8���ZH8��Z�sKX]N��M�]͡�_3��m�auԕ K�rN�"vJ��8s:�:;2d���Mc8z�s�����	A���R�_NX4���F�ZU�||x ��`,�쵔�0�g�a�լ;����������>����h��ĵCD��{�="��I�L�y�� aN-\�-C�d�^$�Rr�ZRҾm��_S+�
~vg�A�����R�$)�´\'[2�T?)"��ČIy �pHE߇� ����V$�� ��@c�Z���љ������h Na��èXk!W�`.��4(] }~��:�譗e@6`��6�`�P?F#�Q+�R���g��S����/�e�-TIʖ�8:����"��¨T�14I;���evW�N������.6< ��X�^�M���0%� 0	H[WB�$)��aA���Y^!Llm��P�:Mn(ԤraI0*��ޱ��l!&�Xk)�j�r�d'{v�hC��@5���*�,z��-2�]iT�N�����ɀ]d�Z���}���Aŵ���p6q�{q��qD���e �u�ϥ�bȳ<��[s2��h&��L=�CC���X�Vh�%�E�������Xmcy5�7���󨷺���Lؽm �vm���8�m}���K��P)FM)�>l��fO�^<x��=��l=��PDv�	RAE����ݬ=Q���`v����(y�`c�����bcA Ȋ5��߆�B�t�ӭ��5��qz,6K��([X��k)lY�ʢ�G�Q�2A�Z���¦�$�����8}�-��4�s��Z]y�� ���Ʃ*�e��9l�:��}�pݵ�"f���B�56���x#*D	�Y�WX�T.��'�]���,��P'*�4�5�I�ku�,�
"��,�TȻ�x��W�G�P%��9�⟌/�m�<~B6i:M\y�����kd
Y�f�p�8�:����."~���Xa�Gg�����$2���H�Ơ�g>ak���Z�O�Ƈ����.�yg� �sL��Rk����-<������3�r��:q�?>1��<��,���g��U@��i4�u):�y�d����A\���h��5M$�A@Wi��ɱq�B�Ԏ�ŵz��CȤ��j��_�"���#��Q��Xt0^C1	�|���Y����P,���{�i���=G[���E�W�%����a9��w��{�G(ל(V�*FixجW�&n|��?�/��o �m���œ/��#3�(V����c�����閐YY���Ŗ�	��=<��Oq�#?ơS�H�:h:�p���Fc�-A���q�0İ�gAPM-���2z�-7_�?�����`��ǿ؄�����O���?{�O�ON�c��(���=���y�x��!lپ]t	.������o�W":8�@8�\��b.��x瞵�r��p�]R%�X]gG�p8Ps9��{�����h{��`yv��|Oj�8�B�Ie ����� ��e���X�C���vb�o�n̜�`n�8V�Qέ��*��VA/'F�ֹ���3��[�J�_�_X�t�Z����"k�����8TOq�`Cl\ ՠ�.�M���	��®��Ǿ�.���$�?�sE,����
�Ocl&)|O[q��L�չ$Q�ݸ|A� �7C���G常���7^;��Z��:�E��Цe.�<���N��=/�u�7m�!h����lɊyt ��r���ͪL�$�ʎ���tȗh712Џ��6���Y-"H�;���O�B���R*� �͗��O���E,3<���-��]�Mbl�YbG��+zC 6Deʭ2p���QTL��t���U�M����T(b =z�N��\(�Y� ̳��*
dCI��dX"Y�"Ѱ������`�.''A*��ٵ���:�I�\�k�JC>�?�����B��L̺Xʗ1���J��J���:�*�嬦E;��p遽�<<��x� ����Xw���u�N��x	�p:Eচ���Z��cs�8|r�J�Gp&|v���Vo��������V�ygQ�	��l*)�8J���6	���a�����.)~�;��.޷�#a_U�좀���~��[-#*��Eh��t�x�Ů�QAJ����~r�_ϗ	N�2!��s��_z-r^,9��QB���p+�܁�4�`��}B��:<�6�v�˄�N"ɻ"���^�G��};7���0���U)� �"z-6h��Y���N�rE�=�<�nD,J턗�ȏ��4%l �+>G�_<�Q?|9]�[Ǧ���iT]��QP���i��=[p`�6$��:��l�)8�߽�ї��� r5���*���M/j����"��N�o2[�eZ-�܍S۾�����=��Ov矟�N��Z6�;�������}��a���t��R��zd�KSkZH8�&�l�����Ss���E2���n�_��̓}�V�x���q��C�<*ȯ �F��L���H����2v�،������ ɘ_g���m�L�8���x����T�6� M�&�O�_�ki�S��.��Nr����s�D�Yv�x�7p���O=+�;_ ��'yks���B��ɪ-�~�-���Ʀ�a�Ir�CاဘB�R����4���?���4u�8U�����l��H�fU�=M09���1�L"��������W�����1JE>Ө�s!A��8<<�͛&P���0��������t �"�XS����|�<˸֦��0>>�I4�G�>ƿӧO#�Ja��͘��4��l�p��ƫ�-�R���P,�qť�`j�b��
N��uB�&d�|��q�7��J�$�E��B�NQ6�<�$��=ૅ6��K��p�u�A����|_�z��UN��x���iD��뿊���Z��{�C����1���J��l�� ��󿉑h��*��=��Z:����'�փ�G��F���j���ۇ` j�UPf�������g�;�li�d�ݷ~����߳����/V<��|��q��p�����xb�?��;��+.��� ����/��R��1I�4��{��?B��$���mINE���g��MW]�}۷	�I�Q�1��`Pq Mg/�����?�R;O�u����x�Q/��l"v��0�v\dnb���s�/�D2C��Z�x� �KY�8���N�i�RSh���:����_F��yM�X�QU��R��chu\� � %b˝�Z���m�p�8�da�'�XꆒQ��[�Ax�Il޾{Ͽ�ѭ��d+-d�U���c;!��9�f���lN�<ة�؍�M�+u�}�j����"� �cm5��_|E�d���`��wk�H�]0�4_f��Ȳ �����}� ���ykB�s�������2�}��(7*(7j*ԡiw�&o�x|�016��Sqժ!@�!�򳅔��/�`v~E8�>�PXxv<BA/��1)L��T��āh4.}z&[<@	=��	sL����W���5G�L�F�����$���}&�$�^���K�d��/R�h)�Ù'\+����4�2�r2�X�9S�C�/����&D�ZC�PB6W��jF�5	j��Ӕ/�sc���H�}�{D���Z3+,�_���B�YG�����.:{.=��?�>����C�F4z*W��4��;�^&n4�|�lI��KY>5��\�	�4�1�̊:�͚��x;�ߘ�ڂ�v�n��	�~�Zv�,l��ڶ<�=	�b�:y�V~��6t6쉀:���[r��&���^�K%t�daG�I�=��Bv�8��y�(X�G�!;��eK5�h����,F��$x&1�t_����e%Gv������!�򺙘�[Cx^��G����p��;6�&\ݦn96s�f96K-��c���4;L@{��K�`��F|!�Ԓ�@JB�Dne��B��M�a��$Ws5��[��sH+��'a�J9���7��K.��PϜ��]��K*ȑ��)+�� �`9��s����çe�F5��Ã��A	�� �^��ɒеȕ�ɯ�$���~h;Y��V�iI��	>�/6d���^���.�8D��>�߆o�
6����F��2�EzB:M1`��Q�!Qb���KDQY[ų���ǎ"�P�ʪ�	l�e�˟R�:ȦB����v�݆/|����k��/&�nrY(.B��&
nN;������D�@��>�a�N B��O	c����p��	W1vBF
Y�@$N��#�.�{����;��������.�E]K	ʚ2RƲ�k��h���]���O`d�DW�Eio�<.!��0��$������E���#J�q5���'m�&�)�y���+V>/�v��S����}=*'z��,2*�1oI$�06>�\��Ϩ�wt[h6*��Ţ�Kϗ�V+F��
���
�s��c�A�����̌�G7mڄ�۷[�3��ţ����QA�{ahpP1/�͊��N� �a���*h��&���	A�y�I<�G%���Q�u�l"�}f&f�c,��%�R��=��_�#��}�"�K���>�;�q��.ܾ�ԉؐk5���GB��-�_���#�o�;�<��_|�up#��������oo�{/؃�׉&���T����퇾gdŶGfVQo��'�׺T�#���G�pHk�0v� �U�m�}w�r�_��߿���~���+�z;��C���?��p�?�srvo�u���GP"NDB
����	|�;╓+��IHO�!�/W���Ӊ���ƫ���Јa[3������s:m4�)�F��i<��)�U�pc���pQ��x�-�sH������c0��@�8�A�&��k�V�rN��x�簶� 8D�A]gKw_̋ZfK�'Q\Y~�h�R.y���f����C�6����JΙҼ���$L �׭�q�JB�ny%C�;p�ڼ����۲K���J�fӘ���V��t?Y��c\��3�{r��^���$o��XZX��'P��st�Z�G�������I�� j�V�f�ϟ�P��c8:'7Ȏ�B��zl�$��q�5�ƻ.��R�@�x-�V��v�&'é�aL�Hn��4�5���9N��[���
��>���Q7r�~���	�$	2Y�^���	ǌ�!���5�ă�C)�,,.c���N[��M��زy�T��)��!Y�$�T=`�Rl28;@�`�Akj5�T:�r�&a����aL�� �:��H^���e'�����A8[b�i|���\��T&�͏�'N�¢���*UM����6#��DGdf��R��i�^\U��%���V�������dOa�� b~���R[Q'�J	]��s����ۥ���,����V׉\���tY�Ǆ.[�[��.C �,�������̬Cg,����K��V�hC8d�g%r\��S�z7�"!���1Q�ђ~t9�p�{���V2\�.S�>���2�ki�([+�Ɇ��J�-)[�GΨ1�\��B������wE	��`"���i��2dlө6ɨe<�5)��mQ� �q46��V1&�^��y$��#g����@{��a�Y����ER=U�����S5�t��d	y7�����r�:f��d�-�Xׁd�}	$�~��E	y�m��K��|Nĳ�j���)<>����*��$��+�#`A05֧��G�I��Є�G1�2�U�+=<��WWQM�2y��ĵ^d���nْf!�� �z� �ɾ�^�g����!��	���ɑb�b��^������x8L�YXҘ��j]ym�z��QK�Hs�Рr��t��"A�3kx�'?���|*EP&����_��̧"[�q�����O7��^D࣬ ��e�Ra�F	��l�0[�!䇞9��`&��flI�z��8�!ω��0�&�T��}OV�J��r������/�/��-��5��T�Qj�$\Wl5����������P\���o4���ę������P�e��S���Ԥ�"/s�1G�)�Mq&$f�1p,5 �$ľK�9����pziw��}�y��H�e��yo
F­�R��K�P��Tp���'e�rAf���I�[u!��UB|H 6S6�Q�����#��kl����YN��F�a�DaieU1���[N���L����)�<u\ӌ��1�#K����8:>�`$���XYˢPi�����p��-�~��nL|�!�=��/ܿ���_v �v���x���cf.�B���I�(W2��������o����u����������r�!��� ;7\��~�ո�}��^�������~�����n�Z��׏�"_j �������`*RɲQLwO}��^��T����]?���{��O���tջq����6:ddń0�M��7��_��}�t�#pGcp�����w�1�a��8���.�ܼ]��¢�F�G�=���n�����'�;����� 1r2d�_����V0>֏=gM!A-t�� �&yTJ�zp��	,LϚ]�������DP9#� �ת�S/bm�8��54����U��!U�TB�x�($.V=d�9`'�r_��5
f'�����\n�p��Í�b�O!���|�&�6n4��[w��w_���Jm O�F�!�>%�L	8�cd���m%~@i��8t'���`&aT�;r�tNZ�RBm��!�@wR����c���0��ˆ	�!?+eGd�(�(�[7��T���o��E�g_z!��)��פ=-R%�9�61�L`����c���c��`#ф8#o>�16�B���:���GG��irL�b�)���4���W�A
L���g�|�KKH�
r�dL��XT�"!8��y]�&��Hp��I����`�b�}���[X���'%e:9�	S�&ї��p�$~Fve簖��    IDATN�ް��nM��+˩X�4JV���'N
�ȃ����տ���C,2]m��\8������I9èy:�	pٹga�н�t��à�TW�z���ujϭ�V{�+f,��P�
1�i0�r8QhtdV6��aa%�b�aГ2��!Ɓ����"%^
�����n�U��� 8�x�硱��$UNd����mR3sg��_l��q���:P+R��"�[G����֖TP�4�� �% :SZŃ����T'��?$�?^wWe���3W��:��<$H�0��a��D���:�5�P'�·[\��\{�ᤫ�D�A�����^�P��lՐ�15ڇ�ݍ�c�����$a׍?J��"L�h�������������YzRT4��U)��E"�TA�}�(6Oc�?J�\8:�D���)ȇ�B��A��������C&_�\4��#}1\y�~��mɦ��MaF1N=�99=��χr��L��S�%�|�(N���A�Ѱ�,��$��Lf����n[�'�3*Y�����҄�eȾ�3^vqa�+a|uk�d�3S�s3��޵aEvajs(騉c���)kY~5���0M9�~�HI�F�f��\�
^~�i�>x�n[>�;�5���Mڷ�L�wu�m���o�l�u�\������Z�&,9;��;6Z��<q�L�L�C�5�N����C�H�g��s��H���Hؤ�V#�1جw���M���c�q�������Ln_N�W>@�����X@6�ZV���7	2491�zW���D�%�/�y�˰�n��H��b�qL���	�Y)����R���+��� ���{�h�,g
����qǝ�bzvE(	[�����-yѐ�luv�{-q�&ƇQ';������`2o��L��sB��~�TY�Ĳ��ӧgԼbG��!+�]��H������U����W^yy}�&���V�T1#O �!��ˏ����L�2'܋9��\Z-L�����p��{p٥099�`Љ�t/��&^|�~��A,.��X��6�%8�e|��_�_��籜i��'��#/qBЃX��:VgN P���\�����8o�4�@6���ދ�|�[��r���Gg�&�rDrj]���T�3�VuHƹ�Y-��:��_�������4���_lB�L�������|�>��_v�>��� ���=��)��?|/��&���yѮ�Ь�0����_�����"�'|��N.�������4��ޣgA�YÓ/�ZэH��Tb�6ҹ��y��$!���+�aח�YbT�}�ſ�ӗ1?=O��dЯ侜YA���`2����ԅ�O��I�Yʓy���m�C��׋-[�h"@M��`2�]� R��-�T"�!�\��IXl�e6e��M d��BȪ�hE	ǆF��[0�u&��w,��BQ�L �<���C�b+�5�R8��@� QrO�IV�ȡc�k�x#��(-�D��L��a.Vv����V�eT,25�"U�����r��d����X�;�J��o�.��l��.����y��{���j�U�`jr��٩�4�j�]0��Ǐ�B�م��Sp�{��FU���Q,��c�!!دB�Tj��#1��i'M�� g�wi�477���j��rrdE��PJ�+�.�+h2���r��U௔� ��Ѝ��E�r����!L�����֌y4v�]X��Ҋ����pTk�I�@��"%�J�2V��p��G�z���`C#I��T�6=�DU��^�St�[E��A���E���������A������L5:dwGD>vlVBv�F��q��]Ҁ�&���i9,���8$y��SR�i�XL�U��E�v�u�[��3��R��zւ�
U78�z������#l�1�z�N��Q�&��yx��>Ƅ�P�B�(O	��[/O�����fv�+USk� �0ԁȢ��"V�2�i$�BW]�7�0	��j(�}� ���!��c��c{�F%��[?�a��@,�m�a�&��M����n�bQ��VA"Bdf6���5���<�4ڏ-�Cr-�!�g"Ԃ�����vWI�׸\%�(���xGO���4]�ˈD�	�Ѭ5$�@���[6	81����U9���I(%�]���XhJ0=�مU�,�B>�n��vMat8�(9L�(�H�{��"øD�P�6Pn'�s8��šC'�Q��� �_q^�/!����NXR&6� wҮT�ΞxY��S/GWE�q:>�b�n��;�51�gT�X4
��uH�Q��J2M���ф��)[V�� �PY�.��O]ɱ[&|ƣ��lN6�ig�ˉP�ɜ��O?��o��^��F�Q$�۪Sp@u�9�04��b���}|�un$�)�p�X���0vi�����9���%e)�pX�"����.�,OM�|4�
c|xHg+aH�v.S��	_G����b'O����
�
�tz���E�L��f#�͙6�.Ɵar�(�}�e��s�&	7��$4��dV��i�̵L�)7\/N�wZýJ[8�1��?2~F<��;$��aH/�GI/�h\~�hp9p��|�λ��%j�x�p3VX���3'��*��H���c2�� �K#���^��I��8�|}�3�+P*Y�$[+d(�R9dÌ��?�gP3Sw�c>g���pD���"��ge2�'�T;M�q�d�*b56�V،u ��JX�L�6�yghrid��څ�������aDj(���{����w,��P�wQ�2U~g7�W���y���}O>��^{'�id��\^tȟ[]�z����>v�� �Nd�{��R:x������J�FK��=N�|~x}!�!�k�wM�;T3K�s����}ꆿ���H�������o��/:�O���&v��H�����Rx���ջ��g_~=o������p5�v���ބ��=���_N���(c�}9^o����q �p���^z{�J�"��ڬ�֪��k��� cx$��d�	.��%�"���2����'�x괔�:�,�H9e(������N�:��Z
n�kF��z��I�R�:Kč��t4��*T����ꓚ�z�׼.:ҩ�V�ݪ(����\�ǰv�γ4&i7{�V�����o��QL�}�cSh�|"i�[�!þ֖̪�rґ��-3�w�[���7�M��t��:6�J���ë� 7{�|�Lhr@_�2j� S�`��1�m���L�k0�H���8�a����п}3��е�z�^���pX���f:��Y[�ԡ�~r_�Қ�����3;��F¡Qr�m�l� ���~���h�@�C!].k�Lc�"�A8�� �j���N��j �Z�u<_k��ID�w��y5	��J/���ԍx(1���$�y1�i�H�@��v�mp��Z.�X�x�A~Ƕ�j�sH�s�f�p��ך8
L��x�E��\W� B������B���a�Ƥ�Āۤf�/���<fWH�Π�ȣ�_�x?�s����V���Sc��$D,�8P麂He*x��I�8���l��8p��ضiD�0&����^�VSң��q��<r9�.ٸw�F��`�i����Q�zgA`:���>5���-2�!c�DɆ�,�*	�<��A/7d#WHI;xz]Bk5�\����0�i@��]���\���gL��1C8U�$��4��xKՊ���<+S��Ũ�{���y}9�#Q��(���PT�Hb�0�69x�m�!�=��ZJM*�7p�c�"C��j7���;X���h
��+��x�:=��������\>�^ZƉ�e�Y��J^�@\1�\vc��崽ur�� ��)�S������*c-�1���ť4*5I`����sv�=[�~�l^�:��,�Y'�sR��n�NŦo�Ǔϼ���B�axLb���B�K�'��2�({�<��O���!�����DɾR��Z�lb�u��!�T�� �"	�R@��Ʒ�6֡���Ǳ
�@.�@�&�>�	�^NBioEWtv��J�8!h7JH�<�Є韟����|V ڄ�PA�r�T�!_�q�"�iٖ�P��&Z��<�������$�%����Ntju� �5�-�F�һ�̿�b\�CA��5���J��k��<ë�|��#�i�C����Q�	J S�lP��(���_O�G�S�Uh�����D.�yD(*8��K����|��{����d�d\�]{Z�#6\�z���|LuyV8��Y��g�Uʈ�?|�0N�,"F���j�h�"�ÿ�6%P���pt��\�|�w�`מ\�7�/���4�YE'�,�lNxx�

6u�ߚgmO���@_��)�mPy�t�/�H,�uO�(��4+�E�g����������h˫��f�BQƢ�� >x�5��Gn��][��p{<��!����+(V��7q��C[6��7܈^Џ�U�ʤ����Ϯ>�K�;�Rgm݌�}�j\�k/N�:����<�9pz��khtz�R�>��E��]�d�b���-�P8{��?����������/MA�������������n�W��������G��˯�C�=��<���$���-/��CH�:�59�߻�V����XY&63,<58g�R���A��E�L�Zxk:���*ܡ�T h@VmT�����8�H`|b��R���.��?��'�dfmq����o�IY'�C�#p�,�8w44)�XɐcI�$����I��L�HX���^7;��b)�h8~ukY�͎%-mp��VS�h��cϘ<��׭�����&���'�r�Z�M8���/�Y�_�Zϧ�n�C,85�=�r�2��خ���h�����t_ؽ���pa��<
�<����(/�@��6ŀ�����Ј�$cg&g
#�0j�[���]����l��4�{|�L�٩���j"�HhĘM��7�`bx�F�=��%�J��r�D�
f�5�&��]ܠј�qDc!��9�g�Ǣ�^oK�he9����7v_�NEGN)���j����o���P�'ל��ouսx���h��b� $��atxcc#�Y#mv\�0�!q��YKM(1�)K3�Ti`zf�LQ�>A�=N�LA`�x��Q�����A�W0)�K�İk�݆�=\�,�aa����j�4B^��,\�/&�C@��%���O��f�P'O���^�r��l���ؽe
��wF��.������r��8���8rt�3�|t\n�E���{��di���b=ѷ�+��A���3X;��cc�y9M,�>8	��B�����k3��VJȮ�Q��Q.�(�.��*�RR�A��B�� ��C�ZG6���Ґ��2�ǎa.W��gA�1 ��>\�0|����(��	��h����u\5_�ŨMb�I�6�JŎ�d�sf����̖��'/AMv�Y�6j(���훰oפ
��g�&(��KU"k*�����l��(��XX+���"N�,˃��R	�׆�K��h��6�ɑ>��m��qjK�|���.3Ki�
M�d���O!�/!"$����={���+�G�׆��iu��-�'��׭���6�D�Bx��i<���XZ-"ѷ	�@��1v�t���h�E�Dx�(�*e�(�Qc�/Y�X�"��4'�$^�C��b�!���۱ԙ�l�W2֞0Dz�����Қ�D�]��'�<$��}�iZ�8��N���p G�?�N��:����
^G�P��U0�l1N������������5�?\n5H3)�Y��d�m�Yn!*t9�ܨ���F�G��m��~�S�X�~f"�6	�\�[RDb�E$!�)6M�����l��E�YM�`�c�bm�&�v�v�����0Me<#�)��lT�e	R�S~aA��Ӯ��W3 #��n�.�u�$::t^(�y���4��
��4�:$��q�ё��56�b�0\>69��O�|9�I����Ԭ&���S��5i��W3S��iҙi%L�9a7^|��'\8�agf!���x���@����9!qE��R��8��d�'�)�j%L��⒋`��ޅ��>��_'O��G�?��՜x�$-�Li�j��H4��@?\�It"!)�l˷�SF
)��4
9����;%�==?g��.7��
�
�2k�+/�ӿ;�:�H��^�D���jf!ζѯ�����_����Ǟ�����Ϳ�;�W_v�徫�{%�nǫ/��~�
^x�f�3�b&����8��W_��wmC���+�}�(��66o�"3&��2��ܖ��r��bׇTՋC'���U�PΓ��b9���*)nD�b�C�������wF�CO �Z�F�T
���2���{����6h�2(�R(�����N��t�h_X�p�Lz��Z�j�x^�/��Y$ͱ~Ќ���k)�r!��H�)�yq3���kb�S�-�	_*��G�\�I� ��v`�������\�5v�}�_�����j�4�����8j/��AX��+Ȯf��Z��<EB�(��r�%�[CD�@���,�)n�L��?7!�
/;i�&�<���]�n�$�,�9!�Y	ݤ�68���@	v1(�֪�UA�=,�d�x�a'�HĂ��!"�$:<:]��e��%��lA�";f��:\���ԫe�4	�bj�8�<����X��g���0��f>�2��4t���>�k�#4J<$�0�m-s���{Ȯ;�|	��(W
�.�'��	#�i�ۂ�3�3X|����v411�ĶM��y����jˉ��˘]Jcyu�V{wnŕ��-cIx�jW�#'�K#nJW���B8t�4�� J�ʀM7�Zu�&���}rL{��&���W�K*���t�|��#H�*pQ���n�!ȓ(�1q:#�h�Nl��ܚ��Rܱd?�} ���v6�{�"0�L�,�0X�`�&��"2˫H--�Ʊ�mt%D��6�y}��'F�'^��T�i�K� �R��Z'��k&�*��7"���Abx�xL�a,�@83dw�n�\!�R����Wb~&���g�l�Iv����'��,�	�T�j�QΧ��l���{�aj,7����Q��nBi�E�K��Pd�����E>v
K�Yt�4SJm�	�Xp��:���>Mp��
���	�<�˂�Eh��F�XÉ�,.�
B�W.�1<ŵW]&ߌa��|l��!7�C��6���͞GO.�g_�j��x�$-�t��脝o���M�XU�G�3��MI� kơؘ�� ���5�Ƃ�E}�>!�bP�M��F0B0#)Y���M5�#��m���c��[L���p�p�:��zx�D
Ut�g]�k�H2�P����~3�D�\Q�(���2��zfB`e�s[��ru��U&��
M����7n��C��H0��QecM�4���4)ƅB����w&�$��9���xI�\�g�&72S3��	��$N4Fq! �<���s�󔿊ϧ�.��œ=�/�F�o�i'���r��4΢[��-���T���6�=G:����9ْbԵ�}��̻<.xk�D^�i-@S@^�8{����}��BQ6Ձ���^�s���Y�^_ιs���%�$$H2�L*��s�����Vmm��Z�\��1�	#�H"�(����FI�C�t�_9ǭ�z�wf|��?�*��L���y�羯�
U�*ZkTAb��4L��k ��꺷&SdM�X[[�ԑ�ݤ�͋h]^�>�믿�R���c�qEg�P����oWt�V]�_lڸ{U+NW��[4�V��?��]ݸ[z.N�i���^F��9L�oqy�jU2e�	g�ZMt$���"<<�2)��~��#��)X����&�����=���b�TjuTic&��O@�>��P�����'�j�:u�2K�}SC}�����~�(C�������/_Ng�w:t �D�{����x
5�p���͠Y��S�P"��o�����"E��j��t��t#C�8������>�    IDAT����]<�����^lT�ߝ�ᵳ�h:�Fc�W��oJ��#K8y=Z�~�;б��1�]����zn��4�;w��E8�e�rk���Ѩl�^�K�ʃ����lv�SP�U��b�X��9�y�R�1�����l��i��Η�Xp^�pďd"��(&��~�;�M�կ��?��ǸtnF�`�MD�r�����Y��+܃���p���@09�����hs|�����M�%^n�1�����ʗW��tc-���]i�Ө��9/�IZ�Y�7D���KCS0���� 3�	۔!�ؔ!~�o;�7~�^�G�����a=5G��Jtujjؘ�%����
.�.!���Gd��wW��=� $@ۿ(z������g��U@ԽRmaiuS>��Ey9ei	�b�j�L�E<B*��0�M��L�Pgspya��G�l7��Q ���'��}�.(Њ�w:vԉ�x%ТO�ym~U����Ng�j;��0�AE�5 �Tt �~���*�H���R$�]� �q�M������VWcS6Dk� n<���N�'L�W�f��m�AuQx#q�gN��A�Յ?A�� �bA?�ڎ��>�3��H}���*�jM'~���pn�kt��8����+{C(�Ud�6�#��C�ᙃ�jCp���>��^�.^GN��!lm�Dg����u[aq3�Z��F��R.�J��=�3�A��}�᥆���;��u��h�K�%�d�&xݸ�(8�B>�E��ޯaп2=�r��xɁ>5,���;���U|*�Xz�ȩ��j�M�����+����S��e�j9����i�d=;:ǡ=۰k�a?�jV�%�Kt�4�e�H���MN�����u����YB�z��П�u(�}+���_ "'�\����Bg/��r� 
�����b�����cj}� ��6�L|f#���$�I�h�L]�7�ұSXZe RJ@��*�,:S���'�UJ�����j�:R`�����֘����Ÿ�v��.�nil�6�=���@��t��]mTXs��cY#[{�fO��0:eQȅ���M
�\\��B�8Q*P*��su0ڗ��QǱ���ʹ��Q{e�Bl�Rd�ز৻���,Xy�-Tj�H�a��}�M��wtQ��s���>�;�׶��}H�_k���dcP�z��Ϣ����<Õ��!�K�_O*�5�t
�9ɣ��5��p�V�$Æ��3�㤛�5r�Rq٢H�b������f�|���"[�!k�a�gM�]�^���Hi��~Z3�.�E��;�?Y�iF��E$	�o1��L*,p*�	T���*�.�8�ڳk'R=	�8�&2�M+;���Ȅg�9��e4���[��rEZ ���צaW̱�a����ѣ8z�z�^xAzi�D34�:
~1���X�ҝ(%a.�{B��W[{�hVdܑ�E��m�N�D5�R�H�K�q����Ґ��n@�"A�?�TBÃ��Ƚ�f��*��i8^Ts�(.���0�;���z�4,�(0̜��ܥ��Ia��s��QC����75���?��߯�����0�_���W�,o�I� �J!_�I�é[8�'�R���q�iIX/�!������߉�}a,/����<�S��ƽ��G�\we���P(V�!��:��=.\^~{bW����$�ڸ:�B�5��kr���[H$��S@F�z6���"6�f�]^��]C�ZP3Pή�QɢU͛�1�N�cn\n4�3�>L)�P�J�;�.РC���Ƀ�� iBSSS��������/�V-�С}�G.��fzG���C���,..ṧ��3O?�'ϠP�H�9?������&��1�>|�ߌR݅�l	]
�N�%��!�)*o��(4�NW��:Dr;�e�H��Q͗��a�[A���� �#z��7W���7����lVr�Prn�S�GW�����~?���tyV�.�&z��U��ѡt�Et9��F�I Xq��63e��Efؘ�X^��"j`;�
�Q�{������D��RNo.E�D��d�fMv�"G��@o����)�4�@�99�ha-�G����5~�mZP����+�Elȹv��!��ȾV��nDJ��q�f�*��(�=�����U�e�Ce��lF�-�ɥ�7D<�4�6�J����u�q�
Ͻ;�px�L�� ���(t}Jĩ���.r�Ƭ��9�I2#�އ���qL�bd��	�ܘ����/#�;����8{aǏ��Z��\�8����1A[�.���e�fTg���u%�kü�	�*Ux�Y�领vš �
��Nt�R�aaf����U�E4+����v2���Q���A���O-���٧ج�U��@�0�Fԝv�>�D��O�S�6�̃3��"[��q(8��:����#��n�ݠ��!��Z���j�X[���������T�EKaC���8�`���l��W!W~W^r�8�>�j^�sǩ	P�̮lH��)�銍�]`�ȡ 5����q<4i񵊬���]J��5�źl�)P�T��)#�[EOO7�x {wmE��D��@��}����%a�֤�_��mV3%�8y��Q��	�����yV�&��J��I�'���\�`7!�xXz+̬Z��C��x���8�b�g;m�g-��@C����`�����;ż�k�Y6f*��³	`6���,��i���ZF������P*�N!�W�y
���<^�j5�����q-��$8��Qa�@p�*S
C��ǣ��R�
xS¶��f����	���bE�/ݟ-s/K��#��K�G�"R�9! ~#�o�iB�:�"��nD�,�Z��:��@��Ԩj���Z�_g�ҍ	k4��3�m�a�`�4�E� �R��&h��t[��������v��k������kh�v3@�� ��i|�|<5V,�%8�|��m��vuj�M���NA/��.���A�>�m�&q��	\�|����μIƓz�l
�6ۺ�y�רյg����v�v"ƿ#����Oׁ>���א�~�\Ƥq�LR���4Dv�18�E�@&_�C�m���|�c�G����d"�:m1�\s�֕M<S_��AFϕz��@?�##p�"����t�IʲO�ג���QC#�C�XhAJ����N� >��.��g�3�E)ߤV�%���?=��O����������/�����.�o��/��%�zŹ�w���rЖψ���"z�^Loŭ������9|�_Av#��~�<��l�Ws?0h3ܪ.֫m�rz��Y@�F05 8$n|M�|F�U��;6򭅶���PM��ӈ8����S'�p�Z��!��Q�o�VJ+���,�>�����-�21���6�*�Խ׵����P�,��A5���H�l`����am�.������s��?E>����_'����	�Umc��"����'���o��d��oL��/�4<�Y]G�e����{=6�U��w���I�eC�'�D��V.c��0A1_���6�@�wq����A�! ����9�M����8	���әD"l��`tvC@Q���n'&������a���ЊPms�*?l
�Iu�(/��\ʙQ���;�W_=#��X|@(+�uD�>�lڍ�>[:)�\����eC7htJ�	y`����%�����N�)Gν�$�R�krQ)f���ΐ&ڋ�AY�T$�嘵V+#�M�T������^9a�q���BX��IP����$���A����"r����?r���U85:�����,�I��VA�Ot�n����%F*B"��hE�\���e�y��F�7�߅��荻�B[�Ѣ����D�]�'Ϯ���0��A�EA&��{��̍�#�J1�n��m�.������CB����\�[B���Ój��\�,�b��}@�IsS	����BJm$�
s���]���v�%�6���Ni5�K3R����B.�x�6WV�~٪�6,=}���>�-�S��g3�RD�qC��f��¦	��2�BemZ�b=���4�<T5]�b����sB�\?z��k:$�I��kj��Ĥ�a����S+A�v��t@E&-��� ��kD����t���r�ڳ}�����ߢ���4�]�?�7dф�>�BE���P��ߥ�b���mB�B~�l��8���c��0M�b�r������,�\E��k�&����M7�C��E��@�`�ǱD�b�H`(Wץ)u���KK8{q�kET[N9���DMe�Ll~���D�8�
K=��M	�%����uަ1���7D٬/�V�17V�! [xC+7�׸�slD屨:L���M��<L3��U��df�h)���4�c,v��{P�X��g�Am}1�_A�\��f���� -��@Bb+<��N��"�7���vC���ǩ�����+-�.r�	���ִ�ʴb�ĽOV������UI�q3A���U����{�Ӵ��O%E�U*9��8���Z�� �� \�y�����Qj�E��笽Hoa�P#��Zt�i�!���f�
/tW��f�d>'M���
��c��1�����0��Ts��~�P��j���B�D�Z��e�ģ�퍊�Ө�D��f����vE����.xf�2ן� �1��`)���P����#���@�
�S�h`fjFǾ�����¼��I�N��F�HCC[�-VQ(���4T�{����YS'f���n��[�A����>�}�4�&x�k՗J!::�V�TV:M�5! H���Y]:PU+�M ̄�6P,�~�@@S���}�p{ec����I�n��[��1�?���?���vg�l
��?��,9�E��zv�_}���]X+�#�;l<��� 6�=��%`:;�1(�eCbڤǉ��w����'�ۿS���>�}�����)�5-vk\M�F���@�z�4^���p�©!r�My󹹹�f�R�/���,70�׃j.�מ{
3'� �E$H�Y]@�\@���L|�Jd�q�zq�-o�G��6�߼�N�8��"�D��=�����-�܂�{�kDix���	�<��ڒJQ�l�7��J9�����?$י���=�wv��`{v��Ėm��x��q|�[��w��O@ǋdr ng͎]g�B��	���w#��ٹe��Ia�+	Q�0�7���A��Z��8�r���kX_�@n5g�d��,PT�qd��e����!�e�)�ݲU���!`iǆ�7c�G�����0�&�0���b�*�6d6n�*z"A�F��0�+e�����d}{�Č<����.��Rq:F�0ЗB������dJ���*
Ŋ���,+Y&�k�Ǣ
t3aHSQ��6��X4��T�X}=18X�UK�0��{�
Z�,�5������6Q
����"a+t���C���z��Q�Ě�Xo��c3���Z�F�T��^��zUkqaK��6�LzS�ni���=;�0:�+�7G&0�g2������e9tvn�`*�¯Uˣ^������>ml/�����o�-�d[�t�F��-�!ҵ�t	ý1���[�/�t����Zi������bu#��t�fqiam�v&�qB1�!��n��Z��Km�
��?��dA���TtV!�f��Q�Z���s2 ��h��:B<�s9��ϡ����hd�lߵ�8��F�J "[, W�&��av�
�T�ψ��D�
Qb�.-���y���u�����-//ayn�h��!	ȩ%�IA�$��6��~�Oi��s�T����K �����\��(R�?��VJ� U�j�}1�?�]��q|R/"@2b�,�~��'��iG�D�dY�p��� _�)Ř�:��F�,/v��!XD���l��5$3��`��X�PQa��pҴ�^B�XE�Q�����@�{��O��8c��m&'-:���)��
Q�403��S��q~n���p���uU�Fp���돨���
��P|N�,�H��
]יG�h���ۥ�iN<׬u6��7�,a�VC����ոџ�%}�M#g�}�8��/Z��և5�j���	q�x�� ŏ�N��9���g�XO#D\�a
Z7S٣�vdp��i����cf�<{�v��Z;l��r�sO�>����S�Cֺ�F�ƞ2Jי���:��˽��=3��u%A�t~�ea��W�K��ψ��'ɞ>x!��Z�
m��c�xf��DA.�e}V�� �J&�s���55�HM�)��V�܋�1Eo��ub�}5�l����g�z�Y{?o�c�N��׎|y�{|}�t8�B��$��a����o�4�7�q��qM�wLOJ&�I���?#c�z�nY.�� P�DE)�s1�����ҙ��5@��iӖv��	h�f{�b5|����@�iP�� b��~~s3#m�����~���ȕj��r�6;:e�aٝ]��o��o��6�Qo�F�~��ؚ0�af�G7A�ق�f�^�>�H4��)�V*q�無�i�{�Q���Q���WE���'j�p�h�!8�{�o?�����nٗ����ҿYC���<?�_��Wg7�$�e�M���9��<�ޕ��@��>^�j�V,���0=���X[����;��c#��*���_V�7�HK����;7Wd_�H���nur�حʞ�+w/9�.���2�!/j�4N��6f/"�i��h"����ʂ
?(l�c.�J�زu����y��������`}3�W����`pp�M��G��F��.,b��� �Ã�MB5�ř�x��_�_�LBݽ�v�mo}��x:�K5�|1�ص['���Ep��,��7_�?<�u������!lsFp���1�� �%���0�3^Ӥ&���!���sM�#�U���p��������@�hS��xR��1�P�k����X]��n%G�߭�@�Y2�ĵmb`�6����`xzs��(��"���c��02k���&b@K�vۅՍ�&�f�^B0�F��!�(>��;ɛxyuU	��rM�4�J.z���Co�nC=Z��M�8�mq�����0Z��P(��:i�ϘNy⺮Ԫ*��YP�AR��A
	7W"�����ur�̃�p�$��T��R�S[B6�r#�������D�V�'O ��F4����3	a�����B�(n�0���gN#O���sl ��6Z5�n�
�İ��ca��_>��T;nxBa�*�;�v��b1Ԯ�Ь������c��-�5��m��2m3���fh�z~v��VQf���-j�,xixe�u
�.�7_��UHQ�%��Q{Re�ė&���Ht7��|D�q8t]s�^�*�*Q�Lce~^闉�al۹��Q�A��植��B[IS��5boŕ�$E��t�S�Yi'm"�U<h�����M�H\��&f3��l������G��m�B؇�A��<r$��f�,��TO�69��d�hc͘��C���k���q�Q5��}�0n8�G� K=�+p�j�+���n�(w�� ũ�edK��x���gS�Ϙ{h��G�T���Դ�v���J5���v�	�`e=�7N�`m�4�Vng^_7�x�I����)��g���}���[@�����5�~j��8}&̨ط���!�l7:J�DjG4�3��+o�F�9h��0�l�,Ꜩ-����u̐G>�lJ͔��i��c9qI�f5�f�ZX3Q�T�1x���x��O�٪ʚ���}c�_�*˫��15Dn�h�lp���v���FD�!��Ǝ�lo7�{wO��'�B�͔]Y�Z��Vn��᜛b�ȯ�~:0�5�s��T�gis����ip�7�Cم6���ܛg�p��E,��kB��x�6���E�-#j���&����&zRq��J�:2:�ϖf!n�[I����5,�����@{P66�^�`�%���^ �i����<`m���bE�
[S6K�p��p��S�y��{���=�܁������a��عc�&q��./.��s    IDAT*_)i������&��>�C�`t|܇lʐ��]3!�����B�eu�i�E���j�l+R��8��{���V�x�mL_�O������!P�~��pS�o&��KN`�,��V��5�f{�,�9�� N��a�Z	bp�a��˥�. 5'պ�Yj6����:���2)J�R2!��7��K��Ԕ0���F9��yp���~�����O<���i���^���׾�������q�ӛB�xS�M��{��`^�oUt�&ǔ�{��yq㾰���v�Mx��a�֭��R�N��[��!����;�҉E�>��P�4�^�TJ;@�8���S�p�T7��nM	ѝ]^����+��3��Kh��(�� �^E�l
�V�HWYB��{��]w݁����Tr����������LLLj�)�M  �3.h!�^��)v�V�@{�D���i|��c/J�C��[n�A��ܴHF����a���Xo�q_�[x�;?D��F49�HlՎ�����;�6n���C�'-��F�����Qt����F$��{��,\�E'����F��)tG�U��]��)�Z����y4)�kg��{��v�!����<J�n눂Æ���ɱ!Ye2,�bF�Q�<�kD\�B�%���M�x��QP�`o
I&n*q��l!+�[&����U��3�6�p'��BE�c���:�ZV�@�I�hժ*��m�5��
C6f�i��Dr�h��hamm�/����bێI��2��4<9.71��A�n��5��AJċ��@'f. W�	�VfC$���>�(ڪ��5��k]�\ǩ�g�}��}8z�D�Hۮ����@.,�w<XM����y�yv�R�`\���DM���LK;Y��K��3����w���i��>	���h#�/ W�b%]��f	���L��RG@Έ��v�JW �뫙��5�j{�7��H�M��_��W� &ǁ�fIt�-xju46��-,aci�f�&�섏:�`Rt
ч�S�0@�!kjF����p�%#$�x�^�^K��k��I�Ԥ<��z	esK�QD��ss�e�2�����|�
��5������Ƴ�5֪OacJa�N�j��3�bSXq"�'�%&�zj�vnCiY�!� 0?���ƶ�|&�4�_�Æ�VG�|���q�yJ[�v6BјV�)�U��:�w�No���\���V�NӞ��,�\ؿ��	�%�
;Em%�R�H�G�*��Z��F������x��e��f�w�%qa����p7��2	 �b���P�Q�If�H���~��p"���ڲ��Z�����,��1���7)0A�gZ�J�`>ZF�k�n�8[h�:ZKR���l&��Bg�[�i�uw�(�.��/���7�ݑ��%�N���� ��\��j[A�۷M����m�"�I�Άў�j��^-��}���h��aq�&����G��j���-��%w%���w=����~�}���܋/ɨ!OJ3�sT����k��W�D�!��3���a�i�9��f��2�Ӧ��qP�����yf�
C~<�R�3K"]��g�TT�Ub>�����I��Ҕ��NKK+8u�����p�i�Apå��S�#��G>���!����!��@*��� �(r�fff��e�<|/��)���>�Mg͉'U��K �E�����l*$W�?Z�R�`�r��х��4�S���	Q�����p�����v;^x�U|�?Ź�9t�L�%_�dvH�+����&
��A���n��&��V��R���q�q���F�6���k=%m��&�ȻR��%k@�oK`���ʪ2�t�Оפ}s�s_Pc��"�rys���~�����+��_=�Ķ/<���E���v��[\������*������	yä�4k5����[�
����ҥE�]>5#�	�t� �q�͘�܂Q|�tnn�u�kz���x����Ө��g+G���P,B�D(~�Iђ�	E���rǞ�g���T[z(�Wp��c�XY�&խ�vn�[�q�߃O}�c���� o��t9��Dbp	�X4���H����4<�)�Z\\�ɤ144��;�%X���}gϞ����=8r�\n�&�1l�gUhLLLa��n���ěg�<���<�:�:�V7+�Dzq�{>�m����F	�ٲ����,��5���aO≔�T.�>���%t��(�a�*C�,��6�Y�57Z^�!�i�p��\�jq�C@��E'�C#���?��lф�\��F���&kT06؋=�[%Xq&�n	� �~=���@�N�@s�������!�Mđ��_Z����e�y�
�-W�H��&g��
N	 v����dum�k�j����ăe��F�./�Yt�8�Ř�BX0RLZ
�b�3U�H�-4inqK�+HD��1�D2�һ�F��Qn�^&Rp��Q��HՕk�=�R��
��D�@�c�z=Ȧ7���,�RG����,��89��ޠ����^�}�Tj]\Z���i�)�?�8�D�s�W9�ff�n]Q���4{�ػ}��BO<,�D´b�Ց˗Plg��87�����C �1��wo�iEK!�lβ��AdL
$
����D��� ��!���ɩE�R�\��u��y��qD�/���!�e�NU��P�~'�N}F�~�4 �>Q��U��;���&�}ΙK��V�yO1�����xuXszIԱY�"�al��z��s�
e$�]�SL���0_�E���hL'����V׈�y����z�]%u�fr�i]ؗL��091
?�:�ذv5ᠠQE"�Q0|j��l7�i�"V`���J�p�v�р���S�Fڊ,<i��\kc#W��r�έcy%��n�K��&'�u4�m�H����	x �����#�Q.glj=^\\������jN&�ӊ�a��Ԙ�Db�I:u\�D�=�i�R-�3$ji�?�
�^����r�+U�Lс[�o>]SX*A�U�vڴ3�56�5�vT�˚Z��=!��d�)Qظ�:j�������7�nр��9���/�x��"u�!#Q�Ȑb1C�*��1��լi���[o�g>�1\d�\�:n^��x�rЙ�5�-$5(�)0���eѬ��**���۲E�"��{��WWã��$6��[`a�������wq��Y��a��������msj��9	fݧ?�q��waj[���%m�ױ�&����^��ѴFv��!���.�H69��=�)&�yZ`����f�Xǽ��CXYY�SO�
?���87��?��'��BF��7=�O~�\�a����ӿ���g����䍔���u�+:8���Ԁ���Ȩ��k��f�_�f�I�_�Sԛ�����럛�\�\i"h��a��m��;w�_����al�v��ǿ�7��]�8=���x�u�1nY�<1�B�<Bw�?k��ɱ�O��k��B�E�J8d5A�4���v�&��׎g?�èTѥ-��	r�$i6�ҟRW�=՘Y$U惡J3�s��6�޻m������|�37����!��?=�7_��&�y��>���Z?���̙3R�c	4:]	&4��0>>����h�z�1�9y�uu�ƃ8|p�~����Y���Rn'���|�"�z�4'������P��r�D|[�=���0h�\E�퇣V������&����PZ_����a��)�|N�v�@�'���t�����u;Jłľ�Xuh��\T)r	+�.���'���о������+#�B�����f��d��ʱ���^��؈��;�ՙ�#W<�c�
p��%,�n`xh���~����x����X\�`3߀˗�F����8t{��8�
U�J%�n�3G��m,��t�xc���6��r:�z&���"����\2Hj[Aj��S})�ǲi�p]�[?b��pV�`2��X��#A����O��k��F9��߃����2�Mnm������7�g�%�b����^Ƶ��H%��I�~��+G�&<��$��I�h������$��g	ʛM�o��g�E���1�
���J���Z��͸Y����fDhĞ֡V�����%5��q��|J�dc!����&s-�  �Uɝrn2����76����l��$jN��z{1<�/�5���U��ƌE�����.��ݎ��~����U�=�YW����'����*^;uAH~�w��d�,bR�8)`�%�r�Q�|nD��">$��łHF��E�ㆩ4�r-��gW��+o`v~�hbѤ	��d�4+L늓������(�7n���9(`4S���>�q�wk�M3Y�����js���D�^E�VF� i�N�a����=�9��O���x��8��#��鹵^H��ƁM���	x��Ѵ�:�E���)�犈����ST+�ʠ�f]v�L�`qށ��O6}�xq
U��ӂ�O��O�a��nK댯��C.��ɟ;|� vl��h��Td�ָf8�,�dY邋���L�)[RWD1d����C� Î�eQM �gf�`�}&-����ׄ��aK+y,/�0���isk8La|4�];Fџp#�n�k3����G���S\��a9]���q��2*-'�
��o���V,?w
�IC�$�'��\.-�8�,�y?T�u4��Ɩ��;g8}}=��������a�{����-PG��W��u��X���g�gR�Lcl7��L�ŏ��Y�["O6�j8]��2ԇ��<~���7x6^�RN���i��,ǵvCNc�r��_ӁO}�#�O��J�!,Y<���I���Q@�y�6?�v^34R���@T7c�ˉݨ����CQ]���]�Xɔ��E���O>���m���px��F8�w�0D)�z5�T��Z5�ٟ}���'0<���6ܤ���TrD��T���hjI������h��W�f5�W��)�7�>��18�Q�Xp���4�x���Շ���^<(�ƹѨ"_؄��҄����(����P����Ə~����+Zσ���I��+6�g(.fC�ό�'O�縦m�֝eMl�O����u�t�c�5���!H&E����O�Ї�����?�(N�����2!�Z�k�ə�S�purl�>$��F�^u�\&>5�8�Cj���0g�j/�.���1��c�t���T��`l����H[�=Lj2� '����;���O>v��&_���ۿ��oyh����g�p����Gy+k�${����������u�͢�|�����3sJ�3A������s�{b(fr:��Q5����	��p�翹�_��M�mك@j@´]oܠ9��[�����<�0�)S�����y��D0rc��i,]8����X]���#�д���wݎ?��}�E�Y��	��0���:�x�˝���+���/|�o���g�	�yX�g���|�@��C��ff]��SS��>=�(o�V4�&U�Q�%[33����Ho�q�[n�mo'��<��o��kobu�����CxZ�'��}�Q��V�:��3dB,=��:`!-m"_�T��V��V����,*�3@5+$�A>��$z�n�ܚm�
=���l��1�5>dC d��P�������0�c��+��
&ɏ��nj�<��"�Ƒ�;�*��ː�^<��,.�c3W���>��'zRI��+I�
S���\�$��	�q�ˆ��UO@�r:��z:����4p���1���yV��5�'�>Ģ��5���^����~RFܘ�<�K�.k���9 �����1>ù�/�7�|DN�6�Y���2^��b�nSEe��ǖ�Q��/p"7�.r�99`��.+cx8�Z�QԘ���
��+	7��&�7������s˘�[B������{%���#��pz�px���T.#	ax�WB�N������>��J����~��1�:sQ_0����u�L5�'���썝h�ȓ�SWh���l�\:���7�k\�հ��@�"��4s%�Mس7�t�.`��C�!�<�y��!W����]
g�.���hW��uoX։:ܩy�M���`ь:&)�_<5ffWo��9!���\��D^�pQ I���xT�A�VʩtJ�4E�lG[,���s�Po[�c+�!l��>C�I57.iVҙ,VWױ��"�����n��@Q��ӌ��ȭ��J!�f���/� �-�l
���)��>R8Nd�֎�����X���3;�%r,�����F�C;�6��XZ,ay%��L+�u]�d*���8��a�xJS� ���.4��>#\�	n��Tj`n5�3������E�X̦�֜�*��N$��̨V�(������	m%x�����eM�9]$�-�V �����#~��'q��,B�B�Q��<Y�G��,
�튣"�Z�vC`'�H�
/5D�M#&��B9Y4�rl�wNmAms?��c�.���}�Vw���ӓ9�#EU�c^	q��:r�5�����?� �{�(��������aSGʅ�K8�Ϲ�َ4j��M�3J��P���}5�-��sM��D5��Ťpx�TikF��U#��c?��}�|ESy�?$!3^
�	�l�/�\,��m���ޅ�>p��F8DK���i��\�;M��U� }.V�ߗ����3N=�Z=�ߍ���e�x�wR��@;݆��ϯ���/����<���sp]������}����S��[E^]^���S<��w$ 6�X Cãz�ex������^���ӧO������\4[��1�#)Df�q�>d7:Ϯ�����8�J%�[�y8<2����߰��a5�<�#��7��7G�M���BGG*�,i�v������|]�\��W&�&�����K�/��8;�2��r�ʖ�R��JU.C���j}�ω�!�$�q���irIH��Ԋ������V.�������{��ɷ�i����۾��w������������;��PƗ��E�򩧕�5��;t�ؽ{
��6�~������u�Q�%S��w������AO�\U�assО�o0��ۋ|ˇ���=~��ić���D
��h���Q'T��.D8R\+(�������(m��+�a��I2����${�����ě޵{&���}" ��R5>��ݡ���(�,$/]��������zFH+Ӂy���
�����'�\�gЮc~�D'��q���	���7j-,�/aeq�3󘻼�#Gn�;�y�F�?�y{�2��h�
7>�� F�����w��V�BQ�:6��9���i�S*�Q��ht��ב�����y���!6��S�i& �xYH&т�͞��}��aű˹���A��pS��9�o'n���cd��W��_l���ҦޭV�(d0�e��|N�4VL��8z��wxQ(\W��/��iCn�
���߫086e� �<���B�:3%x�T��u��٘��������z�u�U�%9��G"�M��g�� O��p��Ff$lW��!&�	A�L�]O�4y{t�*KCȢe9����AT<HX��ц�5z�s�a�Ɛ�����NqzS��^�˃"�K�l�7�Mo`p0�����T�M~�~��-P�����{�/�"[,����E]�B�s��uHcAp�L�����I�����N���BC��5��PؚˋLۉ���������iX@��+�%�/��nt�[���6vp�w���`&"SVc�5ˍ��{Rq2�k(�3@��X0����;v�@��C����&D����֘~��T��Q�k�����j<�\gt�����-�[h��f�ڬG5˾�?O��E���".�=�b��f�z�p�4[���n]�P�X�ɭ��B�%t�����&�bl���t]�h����@�ƉT���L�5pmNnG*dޯ��h,�H؇r!�j���?�T8��\<s]&OFZ2�#�w���F��B��3N2�c��m�Cyz�S[Ӣ���`T���j�/g�d2e�ll��O���Ė�´*j    IDAT�CS�Y�VM�@��
ٰ�.�|V6�u�y�2��
ES�Ky�e����F�06:�h$ �h��<Ξ9'�����1>��
�l��x�hz����gj��v�";�;v
�?�4�e��/Ӵ�kV��v29�(������^�6G��mL�uOX�i��'�Z)(�rj|�r���g�!p�ڨ��Ɖ�M��DUm*��{���׉z%�����s>�G���>���3.�駞E�\7)�.f�0��%��lԩ�26��6z�dҸ������X|U*%Q_���4����T�#m��p�D�Z��\�o_~/�|'Ϟ���G<٣���V[�X7j��>�[�z��Lo�@�^���E4LS��NH�&�,����m�X 4@˿�nR�Ʒ44����7���[�2��h�36��)�ǡ��_�jU�'���c�͋'P.S�@J�5���ކ�����=��S4"���Ǐ����_|M
��a��m:o�_�y
�BS;@���/�ƌ���8�K�}FH߲,g:+cS��׶W�]����Gv8ġ���}���!���ׄ���e�}%Ӛ�ź��i�! ���\A�,ꐱA��ٲ�}ޛ�7]�ܩ:� ������Є�����k�d6uЪ�	�Me�+�qш�w����M�S�gW��zx��������~��`�����\���w1���~�Aw0r�7����;1<��˿{���#x����ˇ��x|A��[������@������%�����F��V|����`*�r�lP�C�(�i�Ɏ���b���<{��mG��6�,v�)�'O�Ⱥx��|n� ��)XL�yk3��_:���E�6� :א��mbh�(��ȇp�}���H�:�b>�qΣ���Y&}�i�Y�^���g���D<�j	�G����(G]!x-$��(��h%.lf�P(䥅�U��>��|��_^\�����W��,b��V|�bpx���w�������
�&J�6j%
���">���)8Ca�u�����V��?��=���\/VP�WP���e4�.�Æ�虜8�M�#����v@�E62�M!g�r11���!���t��S����C{q���E�Ը��|N�����FI�Sv^���uJ.mɑ��h?��D����Zg簑�=sP(�f��W���`ЇP�$r2ԅ7k8A(�����|1���F��9n�q�<l(����@�,y�}��޹�h�������)_�#_丙�1�Չ�� ��Y�u����6��� RL;�dqנ��*���0���ۀ�Z�o4��~�ʴ����fVt=���]�&0���f	�V~ҏ��6e��L���2~���`u3�p*��v��W>�qs�!�#���A8�П����L�bOκ��X<7��C�t7�����v�t��.�p��y�={	�2�7N�YD^3! }Ğ���kt,�ݚ��)S�`B\G<�E[_G~3� �F�����~�ޡ�ט�!;��R�(rl�LH�i�,J����Z>9������R6J��h:���lz-�x�uz|�}pO��I�G��/]B�I��0�&�"�H޲�5�󛇼��n:m��k�e�I-��@ۦ��pJD�\''
,�,��/��M\Y������F�$���hPS6�DX7)(C�p/j���2s|N��ˡ�BJG��E��A� 	A�o6�6�T⡫��-ݻ��8��書<���r�Ed
%�|'�c^���q`�{��j�Q��7�������tQk�Qi���)㵓piqNwP^��3���὘�:(n<��g�����3���?��^��t哟�gqi�2fg/�Y߳k���tO���q��@������8���5��B���׊�	LPO  �5����D�bu�1t}Y	�l�iM	J��ڏ��>SQ?:�,N��C"]��7M �n�ۦ�`�ǩ� "��Ѹ#r�޻o��>rF���>��&���s����/�x~�s>fėlT9b�CWCy�L��I)!�QӢh���U�A4^<{�,����ajj}��W&�L�޲e������B���x���;���h�b*4Z&00T3BMM�T���"���+F���`�GڅD$,
�Xvфö���i��~���+���g4S�I�Sށ��&0�ͤް�<��A�О���_~�a<��+�U;Ңx<N��WJ��2���?��w�P.uv�����W����Z,�����+e�K����5s�
���>����VG$�B�A{`7v�+��%��sp�-��ߧ�ZOOGo����g�e�ʵ&������3��p����%.�������mj�U��� �v0_\QWnY�k
�|�d޾$:�0�td�[E�V
�ǥ{7N�&k�Z5��Z��Z�e�9A����<��W:朤���
h�ӫo9<�~�����o�]�WuWb;�����/��W�<7NOo���p��7����co��?}?}�I4�.����?��n9��ῧ#N�p/J�'�w���m7a0G1�3?�V$)���Á�ۉ�+95K�.������[N���`�S����F���7B5��u̝~��_�UJ#φ�K;1��X�`��m�̧���~'≰B�<ݖ�N�&=��_L^$�j ^��+�Σ���`7m�8�Q'���G~g#@Ȃ߹X������ؓ�:��n�r�lk�k(fJ�Ɲw܍���aaq�~�wx��XI簞+�Tn�\$�����r��FvDbh-��yC�s��f������Ppoہ�F��KH_��6�rF��p��J4�E�Eϰ|�U���ӡB�@� �Z�b�i�1jB`	�<��.�ȳ���p��"9>�| ��ڐ���Dg^��2�؃�-J�&�M�k2�#�s�P�|_���W*�]�)�d�D�P�h�I�!�Rt3���JQ0�S����K�Ɖ-���BUN'D�kB�>>"��P硞���t)D��62��Y�����R.�����_�	���[Z�+\SK�"n���#J�J��47_6\S�[F�X��F/�VKt6�y��{رm� P/��*�C�V�HӁz�%���8��^|n�;w���#��LF�d"��.�Ue���j�;H�jiã=��<J%�<��)x&�J�3��a�ٔsp��<^~��lI���X�JZ��\_�gs�D��6ȿ����"������ΐӌ��U��1���F��سCCC(�Ş�x��rö)@�im�ψ�}ͦ
��6~D�E�*j�N�DꢬyMP��'Ytq��nh�bk#x+Ź����<���bx|�����Y6�M;Aנ�lޘ`N$�^+ �a׎ql���P~�~D>I˴�N�lҰ��q![�b��".��au-�k�i]ۺ�6���W�iU0x���'�a�����pRi�]�h�؆B/kҪ5Q�c��p!	I������π��K�̮aee�R�+���E"�'�g�IVvtʨWr�F�m3p��r�ZF�>� :��(C�N����e���䙳!l�06:(����,!�x���XZ^�p� <�x��Z@&[�������6�];�!c��[H&ӏ�.:��Q� 'N/��Nca9�;�h"%Q�ֲ�M0ދ\ZsnKx���ʂ�nC�����ٍN�kM�(�MN�C^x�uחp�cj8���� R�8�!����p5���ݬ�I���^������?��{�n�E{��c�?����N3ׅH$�R��b�����r:�]��j_Y�	�i��n��&$B"ޫƈ������#��w�n�|��֭��ڶc(����O~�=��\��y��=|����^��g�	�����v�܆��=�DBx���X�����3�BBʭ�$)A�A��I���Ɣ�]�P�pP�H"�&�i�nx}&�altw�~;�^D�G��	�!���SO�N�+���&���NMm����O��w�.G�b>��_�-z�!K(\A�����-���[u�WVW����N뺳��ԚS�f�	�=��ƍ�[�h 3�����GNh�b�%�y�8w84}  �YK��#��#�`��]����9xֲ|���Մ���:<���Ǵ�u{h����چ�j����x�ɳWu�Q�k�ѱ&�T��^ty���L�/�:!��>7��1��hh4�/䮸g�1�%64a�����j~����]Cuen������?x��rǑ�����7����>���_|����}���{��Q|�wcߎmp�O��?<�~����R�1�k'��N����%TJ]��FP����������;�%�앃����7Kx��2������J�I�	�ހ-84�*��s�M�Сgw:��f��E\~�V/#�:��U�7��ti ,�	D�M��=���}عm�v�|N<�H,����6�/�����XKo`׮]�6�]y���A�I8dUXd��4N��~�������4����PC��b����'уÇ�`���**.�.b����6D��0��յ<f���5l�pG���������-W�A�;0�٬Pk���Ku��������l��2��&3!�bT�-.'z	h��5T�*]�6�M��9)����4%N��mzW���<��=�Ć�1;�($�1Q&w�"1���-C����.T���W��b�4;�7��Q�ѥ�E��/�`7�z�h�wj�����I��z����/��j�ShM��Q�6:K� "�Dxɣ�m ���PX�]�4Ʒ�xwr]���L�̰/#�fKʏmG�Ɂ�\����!kH,����>C�D�h�ki����4����B!+��'�������7�(�b�n0�`�r�h0�����щ�����C�B�.�&D���r��uN�7Qz^;:��J��p:,���I�5�S]i����
�܈=~�{���+���_��J�^8�~tQR�09��t�����1��>���n�bn�������Bv3�	A>�����x�Ԕ
�^�\0u��Z����/�-�٢ؓ!E҈���,q!_�Xjj�I�J!��(��e�&���2�g���y�gϞF�RP�50����5q�b�B�]\䴒�Т+V�S����q"@>4Qb�vZ�6'4LE�a����{�(���L�99�:U�rΝsR�Z�-��,�adƀ=���3��26\�}=�Mh	� D�D0`�BK�j��9VWUW�u��Ͻ��������j�^�N��g��{�7<��D2��s��\A,Z�(��
�� ��d&�R9�ρ����c� Z�.X�E�(�)S#MɊ��j@�ZC�f@�\��R8�d:�׃��f��@_-
GF��$;�Bn�W��ci5���%���J�Z��e�u�a��]�A89i�&`�P��"�wrd��nv���j,�KcS�1��T�"���2���}�.�ڶn��ZI� �/����;��u�F4��ڊ������x�R�����^Q��t���TfgN<Mpz̘Y(�g/Ǎ�8=X�4B"�Y���US�I�ͦ5b��ȡ�����i&A�G�/s�G_U9�j&�Z��XF�ۊ|,���_CnuI����{�b��nSb�K\�5QX��x�46L��z�]x�����/�B���#S����O�6%Ґ�DF��%���/S�:�a�c̤K�˭�v�~�p6���~����ʪ�IBO8�^�G4m}N
�+D��R8��%����w�y�Le�]�.�Z�#�ohmE ��}���|��`��U���1LNL �H�5Ѹ�g�N�K���A��^��T�F�<ig�T���`�Y`gV�w��"e��ho	����'{���Vp��y|��?į���y�8���2�����������A�P9#��'��ѣ8{��.����$��bfn�PH����p��!x�~Q�!o�ω��aQ�}�?<�x��}l2�5<'�z�E���L�4���ꁄ�q�#���?��?c���X�$�����;��b	�]�DB�"FnQ�IAԌ��ٕ�k�۽>!P��@:�e�6X(|l���A�lF^��jBM����N���U3 ���P�x����M���d�	;$���&���r��J��жM��ч�|�O���!�o�~u�_��3U�eock���Ň����ك���N͸z�"~��_�ĩ��=ٱ{x���ꗿ�ɉX�sU1�yǑCؽc#���Ԟ��%|�zdy�y=XJ�q~$��7VQ�4��G&�C��.`!�>�͌��V4x�(�R"�R"���f.����%TSk(e��xPE�lV��T2h�@ؼm��O>��턭\���	P]Zi�D�q|��Poz{�d�`�<>>!�OKs+�u��g�ٔ�G���2�#�d�ɚ`��qD�1�#	I����㮻މ�@��r&��p}tB��%�f�pcrc�XY��8�J&?Z��c���p�7�d�!��KB�`Í(��X��`���B-[���I�^�Ģ0VӨ�b0�R0閚Sc42�pM�#��#�v�9����1�"w�\�`d�"];M5�ڊ;y?���R�A�ٛ$~r�iv�~?6��nC.IY�<Hk dD]x�~eVb�`)���4�<u�X,(\��s�G�$[�BD�����}�16q�UjJ����v�	���{�0R�U�@��,r:�p�<����Ȫ�+�4MyB�Z�a�o�s�4�p�*��Ƥ�'�J�Gb�9��3�����L(���
��Q�k,B��h"@�{�,�=����V2 ���ի��󶭛�y�:I�j��\�1�k�C�9�h�V�u�#0�~����w�	1qb@.vŽ��;;�V�Z�ɖ0>1�h<#/��&�#��(��ɎX]Qϝ||<�覭+Nkk��T/�,t®~@�$�T2!X�x4"ϟdY�b���M���Q�E����#G�|�|����t^K���wbu�*���B�M�\o!���q�kſAS��b�b���s9�</<���^q1���..�&�V���S��.ކ"�l�؃��&��Z�(��R	��&&&�����ٍu���W���d	�K�vu�}:v�s�$�"m(�`�^l��P��n�,fجYF&�F�jFd�U�k@�X��"I���nooC���x�6i�3���;��-���gs$�W2NxD�TZ���b��~��\c=B�7W�.�~۝>�54 ����[p�ڄ��c�Id>�®�p��n4���RHg�|}��>��� �ػC�m���_+c|f�G�I�u��]�oC)�AduED%��������q`v��c�����,`"\) �FLxU�B}�
���BA�$�&�%Wܒٛ1+26�jTTc�|LdT��Z�����M���W�Z���.�ղ8��)�͟�)$'V�q	/�RN�j.���߉G?��V�
1m�ri_��?���Q����T%豃^%6��f�d0���Q��v����g��"�sr1�5e����������$��&�+�T6N�z�!���q�����@SS�4Z8��¼XU�"���t�l^��{w˔��������_L���l�-.gxx����>}�s��/Hל�����BH�OOmQu5
<1_�I3������ȇ�k�X5"�,��ً���?�����G��)� (���߉���'�@�D7�*^y�e|��'1::*
�F�E��,hҩ��_��PX���E�H9mX�S�ދ�=4�D����d�aA�����M0���G)���9�^�ի��q��w�/��/008�\����~�x�X�dEL �ɔ��Z�c���HT���H;����)�{�g��ʹ��ȃ����r򍍀�+2�i�|UU%{���T�+�a/U��y�����M!�K����]��we�K�=�*��E�B;6v}���w� ������W�~�4�4��2b�p�ߏmף;`D�\�|ǎÅ6��އ��N�?7&瀚M�}��[ZZ�l����t�պ��Bt-Q�l��L
'�O`9Z�3����ˊ�����ϔ��n���U-�Z]Etqˣ�⌴    IDATW���th�\L�kL̄j4��u��L�ރ�>� ���{���$�i��+M=�D&�+׮�[�='�d�m��H>�NI�����=}�4"���:�-���G7C��%�V�R�D'�Ue�>��BXYɄ����Cp����.�(�u-Ǎ�)$�Y�L6��6:���U)��K��o��w�`� Q� S� ��
�Y�/Nv���m���!_��`nd�XV�`��Q��	��y)OgDv�X.�A��|��$9a4�nC(���U5��B�cqRU�G> o[#f�9!�� `BBK�RQ�:�,u6��Xj�8I4$��r��wd
���n���f���g�3���3���������D��v� @��^+���jMLFUa��@�N	!5�� 7o��l$!#��)m��jH:)VOY�K�B��_���=�
���������N.ﴸ"�`H����zq~F�7���p�L���7����!(t^�R[��ǋd��ɩE�$��Ĩo��=����Z�)�&­��Q�r�t?5����+�i��_e5e��MyP4�Y����$(3�n;�n�L��<
�Pŉ�M֬�PQ�Q�wV=5�RJX�K'��8j�_�w�CNG>/{���Ʉ ���chh���'D��r��S�Ј�Ⓨ��uID5�VI&ד�F��I�-J"\���B���s�H#��ߕ�Z����N�*���n��R�J�J��)�H�!�,Zy،e�t7HA���F���tZ��V191�kWG�ɕD1g`�]=Dp��`s3�8a��D�($p�@U1�;9���ٱ~��z��@	sn3���#Y�X1� �@�J�''q���ilܸ^��8����T
2���9ȖL���;�U>0kQ�7T�D�����ᒂ�X+�鰈0��;�V����Hf�S���XKea�:D]*^���^��]w����|*�l����'q��9t5p��;�n(�t�Y�`rn�^���}�0��C9���Y���`5��m�oCs[ 7�
x��U�N, �����(���"JB�dLyI���&�7j�vs��)��Ĩ֓A�^��v��rv+���rq�X$�x��_!9?���)����2�P(��>6*��S�È<�� >��`��A��,Μ������KW�e�0f1Y�椓됰9~�X�d��mҽ6�H2�)w,Acɼ"ܳ p����	>�7�8�s��I�^�jiD��W�D����N��%5��u`�!P���K�
i��yr
�
��p:��>���ؽ{�\��Ąp)2��?(Ϳ����+W���D$���(��ɳ]�+�9�K�+�����>���`�d@*S�o��w~�#��W�$�3���|�s)���O���x����PTR�/��|�K_�	p�\6��a���^��SA!Js��J<l�h�9��I�&����gB�cc����}�u+l��zA�{��0Ꮿ��Qd���������He�x�?y��դ4��U2	饱 v��A����ӏLN� �R��hD�X/�yC���]� gs3�~�ٚ�uQ�
�T���	79'��r�����g�K1KIx60(�B�'�{���k+;7�|�C���?�]R��s�X��_~�aW{o7`*��`]O��؂#{w �UNo�p��|[��o;�ͭ-B
���0l��-��]�PRf-�2SϘ�e&�*��Ud�L,��ʩ��D��5����z?jƒ@�,��K�w��d$���
⫋�O����Jr��yT�Q�~ld.�����pz���3Ё���8�k
�4�>�t]��B�+�Ï~�c��`۶m�Ŧ��;.p���q$�j\��Gss#��:0�nP�諡�B+R��ˢ�_�-.,`iq�h\
 v'��v;�l����x:�Y���E{{~)�s�KA0zc�T��Uk =�a��È��X�AU�Jg�ҭL���nĝ��6_�����Q^[�ݐ���D�F�C��B�����<��VA�;��4����%$?J���
;:N2�n��iLƅӳk�Ȏ�;�%�,7����''�*�[,h����As��Ax�UuM�E�Y��%*Qհ���̼���H���I��.�H�q�j��@R�XD%Z�i@~�t�D6�A9f
$��vv<	�bW_�
�K��?�κ�4"�t�dڢƋ��J�S����I%��ت("��$iF1*qtwt
ƛ�NvIJ��h��`�X.D��S�9�5}^<n�n����G��m�0��&�#���s`gkݺa�_�M� �8Q���L�x��ͤ>��J�?�� j�ӌ������_3_���Ѯ�&�2��YK�G���y�V����C���Vo������`�@(�����0�Z�a�F�\[T��^�8'�U"!�J�W/�Y(e�5�XI�$LM�O�ߧ_���)n��i��>n����SI�z��`|�Բ���M-���K
�{��\1�VΊw��PZ�vb��t� Sޙ�eq�����{���%P���.]��b�S"�&J�*el�x\f��m�pw<�
|��V�xe�A=�eFg�Fق� �M��7N�f�c��h
`,g��q(o?��*��p�J�J��$�'��Y�b�����&x=N���8!�P6SI����$�&���Kk	\�ō���3�>�v���މ�N�L���N����W�����}X7�֒�Y�O���So�����0��	���T,,I���8�<6nہ��^���^����&�IP��k�p�v�zJ,=��t%����Hɶv��c�4�#�W�6�8��@Uȧ��
��|��ȭ���CO� �ȓ�$�'�͂��Dĕ���(�b,�{`��a��r%�|���FF'��v8���l�������eZKN�����Ę�T�w�܉��6i�,��bt�:f�e@�WG/�Z��s����"��e]5��U� %Mʘ+�P�bg32���o(a��
ZjFC0 �^8�"�B����4�ŷ��<��;v��@߀ȉf2Y)���payyY�t��I9��%��<�U�BnWr�"b�8������᱇އrA�x� ;~G��N�<+Sv�f���N��/c�uR���C�Lǂ����?��P)���DrZ��$��ϋ+;;���ݒ�K}Z�����[�L�'æ����8m�՟t�4�'����06�;��@�>�臥 �3���x����ɧ�������bZN?M�1��7B`}�:����]��o6��	�;��ǇlbSO -��}�75����d3�D(_N�)�%�\�Db(�R2Q�Ϧ&'��A��/pY����&�q$���7�8u#7*����}}��}ב���{�7���?��q����Ó�}#Z6���.x��8]��ہC{�c��A4)SFqAePeuOMiJ�1b�vUL�XHE�J�у�%{��V�[�`�9�LW�0����
�V��p��z��A�-Mhlv�q)�afl#�#������ER\&�Lx�|R�ұ���mN'��*�zP��}{w�=��[֯�j���0��'ß��ghk����%x����&geˇ^�H@�flij������bm�.����fO��
��La~~��>�%�\�~�!��$sy��c��Εqmt'ߺ��˘�ZD�l��ŇΡ��}�;/T��!�) �)�=�b��Ǫ\�Xe)��^�!���E>��ra(&��M�|��Z��*���C5�\��A�H��pz`�AD�5���b2�o�1&�7IA�MC�&��+�?v\�ɤX�����؀vŭfص��j���S��L�H���ǿ�X
˫a�I�H�&e�h�c��ÂO��2ac�\3�b׋�����	�WϏ��$���h�$ҥ��S�ȓ�;�u�4�l�k�"D���/Ө���hp7��f"�͍��F1Oc" n���%�T�ł��c�RN��p;,�nmB_g�$c�J:L��gJ�3vk6'.�����02:!ʺ�M2*�����/�dԣWP�b��UQb�,�Ѥtg9Z>G��I�Y���S�Yk�j��,�Q(gau:WL���N�4Sړ	�U%�#�^��Hp���-AT��u>w=i�JQ�$�"�����]�F9���}�A�*�XJRhr�zA����%�=��1�� ��8�I�TfүQ?4�C�w�œ���*��C'k�V�-?���U�����M��/�p�uV(˛��l\׉��6�����D��jq#+b||sdrLX,����K��,�v��'R	�j�k��D�	%pO:&4�9��D[��X�p�aVWdXaqm`r_�O���ձI���)�ؿW$>�\&�0���1�)�f��MA�r��06	�ޤ���22��t�U�=	�c�0����}&_�P�)6_ʰctz	g.�`~E�x�o����#�c��	B!C��^������wo����au +��\�����eIV��=ر�_5
J�S6�$�P,�l�:�v��Fk8�1h��&*/�}�LQ��6�@�s�΍�.��"I
�W���pg���+�(�4U3ِM�D:�m3�����^�!���a�F^"��i��x�Ĉ�%Z������{�;��>����`xNo�� �8���	��W��G?�|�G�q�����������9��$Dy~&�A�(�╋XX���x�AI����Ec��v�	�ㄅk��	&�4\�=��o���H�`�T�8����'|ʑ�ٗP���2«�Or�}�b󦍈FC8�F����u�����%�ޞ~uͫ�hll~���H�hL�O�A����f0r�J#���L�Y��+��g��c����C9[��(��_{_��7p���f��A"5'���nç>��8x��{�U<�կ��ٳȦ�0[,h��(��3e���ø��z}b�7!nNg<T�S�,��|&M���J�q�f).n��i�I�,$�LOM`qq��_��_"P߄p$�o?��L��4���o�M��`^O���B�1��5�@�uȧ�M��"��P�5������
��s  ��*����꽴��k>M�Mżx��h���K�O��Jk�XGQ�\N}c~��W��-/�X��7������R����/����E��`o�Y#�]N�Nt�{�#�c�P3�f��i�~��#M�Iv:R� �)ae!"�*������9Oť��/��JY1���J�p�Ri$Rq�+9�7�aÖ>��86����q��65��\���$R˓0Ը�I�R�D6�S�)���.%����$R�{��}�#hooG����2=3#݄���e``��꤂f��BO&R�0�DɅ��Dss3::�D堩9��Nk!��	I��/c��$OT]R��!6=������!��K1�N`zn�ύ`lb^������R<#�4t�c��}(��OQȗoUD�X�V��6�	�(W1?:���`I'�4��B&� �C@%-�Cf3;�twUP en��.��h�dC��;qv��8d2P�����~5�b	Ԉ�5[0��*�!���B����
!W�S��ps��u���M�dsk1*�j�YTةgQ��v�LQ�H���)��)Yo�͓��ʝ�A����3A�"n��#�#2)�4��X�f>�THF�6�aM���������LHHٚA9,�XUY�#|3<n;~p9l"�⇄�|� ]�W#Q,�C���ɧ
���@WZ>���)��Y�d�h�B� ,x��u���1>�Ϗ�>lڴYK����&xYMa,&V�b�8N��.*S?���0�S"���*�L
1�Rqم�L��8	4����r(�ePٝ��������]qv���DH�ZH/��I�$R�@Wҡ7<�x��T�D
�|�MMqd���Ϗ�]��!|(��9��i:?A��L��G����[��25���CU���&�R\F$���*1���ˇ`�Id�+1+�4RK��2uRRlXׁu�:���/
���b�ӌ�����	��xvy�(U3�W�9,H��Hgk�;d���Eh6���n�$����4���4kk��~��Har��H�
(,��+8sqo��$r}�wl�ƀfC^��UY���N�A�2'�����|�ӭ�JB�&��J��u#z!�:��u�a;BbU�"�E�Ë��(�^����Y����qx �nGO�G�L|�]ÅKQg�a߮����B8���c��%k���܍���@�[�Q�O��Fo���Lϭ"Y�!���h��_�
��)��?B�y��ę���B$:)~PS2��0�*���S֍�"���\�BV`�TB!�>��b6��g�����J���e4�YXb�c�@�(}U���nkQ��*P��i����XRX��sWp��ψ���,�[Z�W������RB�t�*r�em��x����t8}�mqۍģ�箻������l�������я~$��=���$���$�I�f�)?j�{�`sX�07���l��o��fl|x��8(x/#�čݻw����O���.S1~}��ߕ�G��	Ŕ���ʵtw����]�l�Rxr��[g�g_��k��X���f
y�E�00Ё'{�>���F������s�.�I2+�ӕ��"�߉O|�q�߿SH�4Z�կ��}��v�k�$�G�gVIf�:��^/�˚���a�ҍ̈́(��9��K��O@�Z��kE��7!�V��c���``�G�Ŷ�۱��ɧ� ���p��4��&�k�F^k�R�R5���S"����ޝAq�����f>`����@�a�	�}���ҡy��)��)�B$L�/�+�zY/2)�{"&s�����D���N���rBOc�Jfmn�@��x��������!��^��O���ӡ�aw���Zf�r4Dk�j[;��#��s��tU�y�Qcg���7p��<��>'|�4[���!V��:9��ٴ�M��6�&�k�iL.�I�F��LR\\;�����!$�+�.cfb�Deh
	�w5��K��hne&#��xت�tCs��.x�#\�~�w�y�o? ҍ����я(c5�Ǚ䳂��}Z�����<��ч���$���[�lBOW�@�l�XX:B�Ț!:��&���N����8���XV�*�Vĕwdl
�/�#_��O��"�_�"U���І���x��͏L(�ɱW�x�M�=�Rd�bj�.���Z�$�"�,*Q����V23	NS����KB1�;5Jw�I&>�n��@Ȑ���w
����M��ۂ`vn^:U�ZY�!;�$#�.(Jr��+t��z�h	֣��>�C�޲��t��i���S�]K��;@D�+�XE�Ȍ��2r$1�*	��3a��T�@I�fg�U>Iv��xX�$	SC��k+�n��c7[��eEs%9��Ś�$��$5Ĩ��&Iz~�����Ex�4��]�\�T�dR�T�lV:ۚ����^'�,|N�V�����2)����0�W�8-��V�C�S} (�E��M�=ݦ6Ԇ�9���
A�d4�b$�<��J���_'�]�b&��fZ��
���8幭�����Ĥ�xQ>G���ia�HWS�1�	��ߪ/��.5����/ѓ�=vC�U��V�[ʱ���-�3��	W�$W�|e r�T��,�7IM0���]��p׭�wJ���߄	�Uu��F���E]I��\N�)m"�)e!���j�6���Z*Sa%+� Z�4�91�߂��&�fdk�Ob�֡\�`j"����XY�(7M�e�2�L�g�JS}Ë����J7%dRqx�fl[?�ގ&��@�i��Jq4��ڧ*����f3bi�G�1�ǹ�ゟg���݁��Vt���p�d�=�@"Y@���V(��LF%��ǫ��ب�b��O�M"�;v���UVi8��X�~��Ҹt}\x[$s�l�0�������,��$�før�
�=�c�V4)�XF,[���Wp��b�6bǖ����ˢV�Y֜TS	EҘ\�ڍy$�8�]BM    IDAT�0Z)�L�#-y�r�I9
��*����ݪ l����,��7S���`"�4�t.%M�5��шH��P����+/!��
�6i��r�6���Pn����40�R�!�x[M���#x��?�m[ש"�?������3��g��ć>�>��G��R/�%����Cb�c�zrb�7p��[�|�"ҹ>�����O�:Z��Z�V���/��^@,��{��&L���8	��LS���d���I�Y�3a���$����(��g>�)<��G�v�P*���˿�׾��$�w��R�S��۫�x)gY�	oCrX ���K_|
'��2���E�x����x��G���?��_,�����'��O~������OAh�H���Gp��^|��Gp睻�Hdp�̛x���091.����Q  )@ֿ��cr��?���c!����Vdn���K:DS5'T���d���F���{	$�f�R13K�*��������y�c0���/}�z�D�i���K!tJ�����zgS��	�-�K�y�o!�,bՙ!�F��Y|1܍
.D���VL�/SU��x���ffIG�PNFa����3P�g�1�$��1�&�E^��}R � �B��:���{>����;T�����ߏ>��J���� i*�TJ��-R�Y��c���.�}�\�x	�j{v��Jh_y�)�;Q~�T�����;cxp
i�����X�N+L�6kf2e��5������,2e�C�z������&�>u�r��0������`�T���G1����gQL��\��d�*�;�N&W<̫顙F����÷�Ё}(�3p9�����ի���3O�&!�^�AZ��6����(��j��B�����@�t��Q��`m������GTA���/��%��T��aq�(xaq�3�\ހ��G�Q��[��2��$��&��mD]k7���&�ǒ)��Y��|0Q�����5,^Gfv����"��a4s_P�J���P� ��@MѡYMY���bRV-R���#�Q���#��ӽ{�<� ��XX\{s#Db�U��;V4�'�y��8'A��b�]�A��aag�p-_��4�%��C�hD<�)J(����������t蕻����ٱr�35�.��92V�Lu�u��l����tb����N$�n��+:۪�t+F�	&1�"Qk���I��C2�����$�|�(���j�Tu�'�.��ь��4xB$ʟR��ԍ��$���5Xqq|Y:��BQT��E��3�6��r*Մ��L�����$k�\�v��;1�ó�cg��v$�xv��I�%!R����R��$Q�8i>����ȸL�o%Q��ўUST�F�On�GhE�~ 	wA3y�� �%����4����	8}n)�0@>���H�c��⇒�c�QM*t�J�0�R�
iPS�R��oeQ��a\�L+7Er�d 	�s)�b�����Z�	z� �LJ��[~@8L6��"M�x:� 0Vjp�-���@w3Z��i@&F�UМ�$k��
a~6�|��σ�&�@``-���{����0��WV�8��I�=v�ݶ�*���L!�2�R+���B��U�	�R�B�+�Z��j�X
>����a��"y�$Le3�*ɲ4o�	f�kN�jf��&��:g�A��ɁQ��!
O��_�V�&����_��Ĝ@ٲ��n؀#� 賋�%u�/�-�¥�k��;����ʖ�8w�N����Zv��� n۵�=m���
���b���,�8w������5
���1˒��!*)��X�]Y�U�`�O�x��5l8XlF$S1$3q��ɕM�,Khh{K�Jo����'a$�����J38%#IL���j@�{�FZ�Sµ�C���ģ8�o�d�L���p���p}�4��h�����L�DK��W2�M"��\�g;�@��%�����H�{�{/�˟��:�d]%�i�8~_y�@��Z���Wj��T���X4�HL(%'KN)���b��t����Jgd����9�ݻW&��R'O���'����Il߾]x�����E����P<�섳111��}�Y���)��Q5Y
OG�P������c���=#b�<^>~/��g�pq�f���B�E�wܾ{�Ql�0�����_���2����|a~�{9z�Rr���I��)��:z�87���	x�>y^z��'�z�;�K����,�dƶ�4���f&'�c�n���/زu7^�����~�H$#�sy��J ȧj�*gu6'!$��V�
�ќ4�U#�?�f� �{�+8<~x��a���h�k��>�,�J��j����W���J#Y��>�H�L�lV�/h��?�[�i�7�[M�K�4J���Pw��>x���N��c[����I��]��(�kȗ��X��f��fF:���˂�� ���n�$����ۿ��(�p��d���C��w�%� c�R�N�F� �{&R�XF(U��\c�i,�ʈ��9�v�f� _�b-r�`� r�8�]��ř	��!4�,@:���K0��2!��h.pX��%��j������܉-��1;5���i�w�������҈����{���tTĠ��.Gmbl$�N�9Ew�*1%�R�(���[����$����䏋���<ߗ���L&"���M�|���P�.����q�r$�91�A"���,��Xe�M=�a�>��E3HĳHf����5`����8४N2���iD�gQX^B-A-�TÀ)-ң,�b��7���UH(��	F�Qk�`팊U�8�z� pl0���m߄w|�!�|.��	���9�fAŮnUU��pJ2$um�q�$�Cr�͂&�5��Q��c$݈��3��	Cz�����%�`��Z*��Y:3�Dn�$$�o�T �]�l���y�D�\�:H�s-����ʁ̓KW�aA�u�D�K��$!2�Xt��=�{}�`�n&��Y4�.���'YD#|�Y��q�$�T]��8�g;��(f8���廬���0��^�'R�⺴��]�ʊG��g�C��6x^7'1�mUj,�TrR&ԫZFP��*�4�E�U��f1�q0����3r�W�@T|�	3`�����
._��J�\	�� ��D.�k��%�*t�֭��>!��f��w��u~L����ؘ$�A����F�E������XF�5!?	���aГ0�c&Zͳ��$M?,�^Vk"� ��̥&Jc^�\za�s��p�V����n��	��l�Oe� +#'�=�}�"�uv����WP�|Zby�d@"������V����׃M[��UdKE*%,�$qedc�+�:<����f���я�[�a�#k��jLU�Y�k�Fv�Ua�j,&���ˡF�q���� ����������I�$J���-Nl!r�b>�N%��%#,E��o*�M����`|�l8�	A�i)HN4�D�3U0����D5��%�عu+�q�>)�f5m{��^z�%��1���Ac�W�<B��}	���(���QY5����"����h��	�p �+��K7�!_�?�f�Dk;������%e�:���V�ʤ�e$ɂ�j��jn��bq���YX�5x����#�"�Jh"9�`A >���b�Â�J����%�}�A��;���H6W���������Hz66��Ԁ��.�^'k<���4�>(��	���r��H�dO������������X��/���B��_�?��'���.qTȱ.���<s�7���%RP�����$r��(���/p-楓Rtuw�����7r:쒛HAp����{��|�::��#����Bdry)fX��wv�qh������q��P�nQ�aA��݂?|�1|�#@�P�"2�*��'������W&P(�Y�,�\���A|���Q�����c\�r��:��e�ຽz�\'?���?jڠ����yJ�x^r!�g�p��>_+�q��S�Wb��i��FĘ+��<���D���M����p�{Dh-��_9��(l.��%�Pr��3^R	R��y��'<����M�, p���oE���� �yzXQ���v��0 6��\L'Q)$Q.)�+*c^�K�걛��N�l�kh���@�R@%�6����o}`�O?}���S��������_O²��Ԅ�YL&��~���L,���l6���{�/^���|T0��Y4��}�>ܶs;|8I4dG����i�A��	�\L`t6��ł��>Z�`5H''�M���[6uS��]��Kg_�BS�	K6���8��E��7�`�T��#��@P ɡa7a���رu3V��E���С�ص{����|W6�ء�7�d���~>���2�g��>'tG�4�I!��t=��W�(}��ZX�gu9$h׎ݢ�R�"���c'p���0�=0����#��A�lB2W�b$�ƮA�o���E8�N!��ưP]��v3�n;�6
��'f�� �V�| ��F�A#�b��M̂�Xm�������vjf�W��@
��d���q�R����]�:�t�s�tIEI�0��D�&���4����C��`��uU\�]�smfS�G P'�ⴡg�Y���(�t�I4I��lN �BF,W�S���aI�v�]�v� �q�`0<T�#\)���L"1�L�x(���_��Xt��n�HP�O.��"Q)�8�11ɏ#�%�,ȃ`w���Y��ES��,v�J������؄Z~��M����E��.<3�v���d09�/ٰ��e @�2�b���F�3U�t8�t�4wT�C�j�M��X����	7W��O��TOqK�!�hqu�t�!܁b�[N
~��	D�Yx}A�NK�"�Q�	!�P��֤[����ū��H��>���q��~��v���g��U�^`)��t�nr��4�8d~�I�ӻQ�$A�\�E�t�Y s���,�J����?�E�/��)�+��D�k���I�E:�2ANg�PŧS&4�BNK]m�6���C� FY�l	�3��A$G��Q�?���j*J,�D��\g�\��|
�:̄������{�m�@�O�.Hϥ��F���OL�=�3��Xe����kYL΅D4��a&�=�ص�M�����-SńqIA/v>�Ћ~�
�χ\$��>{Q�8�>�	9G\�*?�Z�lH��*��n`jn�B	[7o���[�s��zʕ*���i!iڻ�n���*�-���z�$^?y-m]h��9g��B������@w;���t�X�"������Q�4�G�L[�x�3�:�\q�Sc����Ҫ}��9�=NPѫZ�Љ��&x�lk� kkaL�c>���%�&��aw��8GwUY�
'DL��me>@j����n��~�|�?<���Q� �?��/�W���C�`�{���ߏ��V9Wɩc�X)�(hJ"<�LJ�I���G�m!��}����?Cog�@C�>s����o��8�e�V����|&�.]���֭���"x"8{�N�<��Z;v���M��at��y,.�cÆ���R��+e�:uO=�N�:��"������4x��(	Gcr��t�a��M�Y>����wp��(�%�L�yru�����x�>t
����������!.\�&'�|�)����m�.ix�u��ˈ�W��l�s�M:��˧ϠopH�<�������E�n5���Ƥ�ω������o'581VE�ݽ���mS�w���آ���j�i�p+N����oC��p՚�tFd�)��u�lZ�A�!�ߌ�5�ݘ��o���M���&b�����:�5�#K`ee&��� \M�8](��Ȗ+�B6��&&��'���Hi�y8m�wC���^��8#�����Z^;����lN�.���
��Ԗ�ݟ}�{~�ٻ�d�.����wS��wN��篿�L�j��l�'���I�X��b��hڐL��m{p��Gp��9}�i����u�M�loŝ�nGO[\v3�4qXa�*WE'�H����lW'c�K#5�dpIA@�aq�#~��~������+W1r��Ut7z`�&�<q	��)Ԩ�c�Tr�Z׌֦V����dri3��;�o��X��ĸ$�w��Nq"��ȏ�C��kmkFWg����"�i����v�qR�����i���XL��(b MV�@ilB�
��vm߅]�v���M
�_�t\��*��V��C�bez8�۾�v`)�A*gD4U@.S��<�&-6�U�k��1D痑^ZDum(D�R(� ��	9Qg�8X�j$��:�]�����q;�YgA@Q`*vX��,�jD;�J����;����G�Ey�ȟA�;�l��ž4�A,�I�0��L��CbJ��}"[�d�N�7���UU��Ē&�����
���+Ja��Q��/	";�<��ꋺ����d4�/Ovcu7G�#��R`�����.3�%Jk���@�F�@��H\=���N�T��Mf��0�#	gs�b\������nd�K�1��9�$��*{W��r�R)r�jE&CGV-���m@b���U9���81�5O�����p(.u�Y����nB:�(���+��e�D��ؔRa�[4�& ��Vp��Y��py�ů������&���֮���$>;~>v��?�������F���nJ�Z�vy�GT�DTV�DDi��(� �����~
��_�$q����ݚ���k�n�^���:��V��^��A<E"�{wg:�Z�2�{�n���p2Wʣ�O"�b�`{�`5�d���I�Ǳ�1�298شe3�&�44��01���ό!� �ƀ�!����ni��MC�mi��Z���"�뀜��481)�J��If�(�������arn�Qd�8,tb�^4x,�
��:d�A�J��!���m�
�Z%���
�;)σ�����XD(ia:�R�\H/Z�L��*2E~6�*nL-����^�lZ�����r;��p��eї߻ewܶS|R��ȕL��{WF��c���Dts������z�]����ND35�X�����1�����b��@k��Zԓ.�J�<:4T�Lo�֘��P��:�7k�67�pS�~���L޸�lZ C��y�e��,\Y((Y�2���]���h��{�a|�Æ��g[_x����~A�\�=�h�lXMoϠ���e��T�;���}�)�(ɥS"Б��ݎw����C_W��}��I)�Z`�:04����~���yG1
���7������k�n��V�?���7���] x���{E��d����J'�+_��l�BgTKe���x�O�T���X���.EC{�2:�c�Y\^�u��ٻo�pΞ����~c�pz`��NƑ��14ԅ?|�q|���%�4����_9&PB�ss����y6q��q��mۄٹI\�rN��Y��y#Jj��wzb����/=N���
J����<xPރ~To�qR��5���).����M�CP��H���E#IF d�fS�C4�@!_E[{/��zē9��/E�ٶ�����Ć�u��=oF�]N(���k��_����9X<�0��}���8|��������b�F8M(�(��"�J����]w@2��\���x4������hn
�I!���	��#��4��f�����#��2:���
O�Q�ҹxlz����>q������T$�������o����/}��o�Kƍ��z�̪+��A�:.�\
�M�X?<(���	����������'1Ms�G��[6��ÇD�i6�=X�z��}=�8��fE�FW��^[ƕ�(R,��`'#���蓴aur�R�ьx4���9��O�i*���S:��k�[G��T�����Jx]~Y�\�R��-��jÎ���a~vZ�-��.�*8u����I	@�䲛��"'%���hkMbnn Ը�uB����+���߹)[�� Z]Z���,B�Q_ZB��uuX�~#vl�%Z�WGn�d�!�7at|��O#����D����<    IDAT�ܴ�k��a�!iW��55%��F��G%�G>�Dry��
��y���!�*qR�a2��H7ْ��@kK2���&d&l�$��CUMjb�n,��m�َw<� �u,���c'#m�N�e(Juꄛe��H�	��("��)�aU;�,��1����]pk�;�4����#$���?t]��nu��ɩ�|�K&�Kͪ\O�T⯺�1Ѻ$z2�]=qf�eW�E&��k�ȣ�M��&vQ�e�seKT�����>��Y���y�R���Z!AOafy�ʕ�\R�3U�l�յ(����SEp�3����,.���pJ7��{�'��-IK��Eau�t�h>���=Q	*� Tn��� ����*P�h�]��tlI{|�ʮ^ܞU�MDi�j�]�c�B��E��B.��>��g1�<�(DF}�t�Xq��].)8bVE��ܳC-
lhhR���ov�4���n��?kdh�P�z�u�/ Gl�2�ѧS�f�N_��� �$��f':ۻ���$Ϛ
N$��J<+��^�����uaˆ~����ͷ�8�d����`�$����05��k��ǫH8͍�`, ౢ=�ǆ�Nt5��m��e1�KgYq���Jԕj���,X�ep���O�a1s&&���mط}:�0����P̪�,8}�T]k�x��eW),{Oa�E٥�T�xn	�S�@��JG&�B�)O3�����5��ӗr�y����؍��)���J"+q��)���6�Z�T�����2���u�$ߕb�Ks�v�
R�U�{h����z�7R8u�:�V�R$��l�PQJq��"!��9.���N�6��&�Z���G�D)��K�}#aU&3(���4+��~��Jg�8��ܼ�>��oN)���[���N�<+N���6W8rh��3����I�}�?�7��.V��u2����@��L<	C�$��V����T��P������H��k�������>��;�h�p���������ŋ�8r�J#1&�w:(��k��*S�|P<��I濳	Z^���E��M�S���s�}�1>�g�}��:)�a��~;,f��o^~�e<��S�Lfy�|_N	�:;TN��$F��ǜ� 44a���9�m��Π��N��L�b����?x��>X���%�*#���y�ΏHA@�L����t��������!2֬ژ<3��W�ɸ�^3��G�ϒ�DP]M�@��䡇�&��~�3;���Zi��G/�>����dG/~��l:��&d���xͦ�Z(
����/	wR���ط/����c��}hj�A�xI�����<0:6���;.|J��K��{��'�����?����#�<l� 
7*�L9�HG��x��;�G�� �2~���ӟ��+x���§>�0Z�}s���X�ʄ��B����2�<s��<-�.J�%�iMn[��W��]?y��aus����
��={b���~�L�b�`�סfQ
�L.�S�9Lvoۄ�>�!�ש(u�ө^�ɿ�؉c���]o6���Eo{'\6���%��-(,H�Lx��x��l�nx��RX���g�ჃR�F�yqt%�+#�C�߆j,����]�����f,�Nɏ&����C�K[{Z����D�\BGg+n߿G�+.]8�K�/`uuN�CF��L��l�B1/���� ��RE�&
����4�W%�c7{ppP>5�~m5$cS�y�=Ĭ��7��=|u�B(Es�|m�ώ �*#Q 
5��Cؾ��e��Z�p�`�7��1��aV�w��=��9s�7f�M@��(V+��c�5�)�)�yM�ww���11�1�^�DT@Q@Pzg�齜^߽���$��~����s]s���|˧�ŋt>�D��-�䎦_�GZ��t��fezQ`� ӫ� H���E
�B�\op����\�jѱ��T�FQ��O��\(7����`��8��ᭈ����=���$[�
�$i�R�g��*����|a"`W��u��y/�$u �9W�G0v[���$�Х��d�ϧ	+u k1�شu�I���v�CJdv�17'h	�7�{�^�[��"<��6�.�Lz��U�:�Ҍ��.u�V��c@����֩Md`(!�7�5r��&�~d3q�5fM����R��.��\ �Kt�t

�����t���\����\Y�ѯA]C��ג/$L��J-Z:P�}�\�y���b(Jb�ۜ���Ak]�=�й�p�+��fUi�s!_�2�� q�@W� Z;��s�A�u���	��+�0�.K�Z�����݉�:�gc�7%8.ڎ5���]�s4��&��_��r��#�
?��T�%��|�"A�����
��`�bÈ��X�Fɀ�����J�D�t�x�Dh���l�!n�x�6ـ'�ƺzT�W(�Kfb"�˞�8<vo�)u�؈i'����zHKU, �0�i�%�'�<a0$�m"]��mؾ�	mm����EA�*��Tct]9�"{�tj�1�dB��'�L�~C���ۍ��4v�>�]�����5��][V��N���'��;���DN�	 �j�߼,��0l��N]@9iS��T�͹ynm�\�ةS��D4|��6�Y��$v��4	s��D]enG�x�$��F�u����?�e�Ł�G1�|�2c<�4r���9®ql�SF�@eU�L�z��΃ز� ���9���@���O�ĩ�%�T�}����C�" {��a�@r+Ut��EK�Q$�QIZV����I`˺u�;v4�Б�db�+/�D\&���S�E��&f8����ÙsN�������6�xk1�����(b܄�8�$$3Yu��4���0�����U��t�x�a?��v\s�%z��ظy}�����2�cR��p�5W��K/�����K���?��R<����oo��6x�>�����/����p�5��x�� v�G��#?�1,X E�t2�e˖�OO=��7J�K*>U����|�&r2�7Я�����Ĕi��}�װn��pKPR^�U²1�Y���7\~��O꽽�x�õx�/oc�'[���=F"5��"\�'tc��E.��~��z�1,�0�hko5\(KZ�S��1�}O�~��ș<묳0f�|��g�r�J�1��R�B�1�2�U�_�-�`�44�3�8��ᷱ �9�vQ��.�Q���{.n��Vuw�g�%[�`8(�f0��`0�ؾK�.úu�Ȼ"����+���c���Б.,|�m�ٰ��<�$t��������.�O~t���n��/���{�����ŷ�v��
�B�Yr�ƺ�|�������_`���q��N��m�'�ix���^��.3������XB��?�{γ��x2�NpV�b�倏��
Y��N�?o���<D�h=rjkQS���^�ڻ�����"b�$|� jʫ1n�8=$:.�T��������V����M��;��F��v���K	�7�iW2�q:P	���G���|��/�d�14�ڂL�!�"ʎ:h��r u��|4��NdVV��oP��|g̨��0q,F6Ԫ��*�G����[��-9�(R
��#)�P�'a�ԥNK�[�ߑ�@%
�H,fRB>_�P3HĢP;��}n:t�t��v�:o�ZП|��7lG31߱<vjA�/����8㼋�F�7��@4��aFޏZ&�!!�g��jjF����v4�(7�B������!("\�@�=!��X�lĽ2D�c���2K�u��/0Q �?C��^&�>�z-�5J�H�R�M��8)�X����dF�*�q�%N�/��U.2A�$ٵ'e$+Kը\&�"b���2q"f�<��w����ު*�����9�܈s9%w�(d6O���]:�T�M�"I�,>�Q�a�c��.`���c�MU�Fq��Q�u���@�x����9�w2YJ�L��֖"9��~�
��TT�,@�!Ǭ^N�؀j��К�(��i9<��8�30dK�YX�X]��_8NH�&T��1;�d� 3(q(�7�\,��� �1q�3ƢHgG�:rL�i�N�b.YEe@�{��R4���H�L�$��W�ΊH��y΁�(��&���A�-*uP�TJ�c'6��S�g��o����6tmQ���_E�	⡋�*a����s\�Q�	���E^��_���ء���q�v��4��Y�U�>���������GRw:��I1׶�z(�.�3q%w�s�j�y�21xYU�G�V����%$V�	�
R�"'ճ���aAN�������%��חBM�(�Y5��",חQ]����\n�CJ]�x����X2��Ã��!�>x����g�xs��2!<��=c*B�F�Ѩ���8���t�l���L���K�X+X��`�Ɲ����s��H�qʘ
z�"�v�Q�q�m�"����`޹s0a�з(���Օ]�t� �C1������f�g�'1��1�Ա2MerN9a�s$I[�&vJ��2ز���9���#����	�v�dD&/*�~�~�֍��5��}!��7�s�aw���^89:���H���ի1�|L�h"�s�"�_��NnV�UXrt���r��?�^�~�t������S/b ��/�x��)�>�ƴ7;΀��\�D
ϐ�~��)�f�=*�F���}�߄;n�I�i���ٍ�=�8�Y���p�ӧO�5W_)u��-ë�.DIq1~��7JJK�ǟ�����5N��_�[6}���G�妛�����?�0��.��\;�o�~�Y%)*�x�����ʐm��N-yJ�H��!�_%���p:X������s|�H2� �)�F���݉��_�b�2�������E��H.�]u��j�1y�D���n�X���\>�ѣ�h��r��~輸���u��y�X��F���,����w�w���E��e��9���8BQX*O���jOe� �I�!I�k�r���е�uc��x�Gp��sU�!��϶��ہ��J"a%`#Ga��PQ����;���/a�*&\wõ��k�b��jm���z�����t�^�±�^uؐ�Ó��K��_�_�탵�����`���[�ݯ�����$:{z���k�e윳h�0{IMm�޿�%�%���5��wp(��ӳg⨺���w.���)ƍ���K���,|k�_d�#F�a\{�,B�"ԕ�p��q�Eg"pc��!�?�3�����*�2Tx``�'SR�8��e%���n�\4|~�iII��z���ջ���f�ODq��u���E�U	qU������O��D?{Z�G
}M�qt�f��� B�D�>%'	?�GPY^	���r^Iq2K�>c*Ə������P	#�R�p��wD&bfzƙ�c(��"1�|�S�L|H�%�6� &�ڋ��}�Ed�	��!�D�pw:P^Vf*�4���W�ISNA�P6���k6c �CK[?>�b/�i/������Wq����s�I.����@\-e�X�*�f�{�=MMH���(7g�_vB &y:�Qe�ݖ�������Q(�&#:���9����7]}]D�$�ǉ	�OǼ[�A��ݽ=����j2��
���S����Y����[4�!U�YэU3�F2��	cF���]�8r��?��e�B^,B�-%Kx�ԂU��hr�����!gGBH!C��Tt��8h��@2���Γ�g�<�;�diΠ�����vttu6����\yZ$F,1����`D�U*=��Q�r��[h.>W6��U%a��B2u����LZ2��bȩ�{ &�&%� ��Ta�G(EA���)B�@G���I�aV�����/XQ*���k%���B�4K�N�3�y0�crH�ʌ�P$JݕJ�L�e��ބ#�*�����%y�����qs��o}$�5Sw������U�;-3��\���n�O\(*ѯ��g9�Z�Xv���d j' ��Z���$c��'�j��7�.�������=Nҹ������*kQL����	d�rHfd��rr���lg
~���2�Gף����2��f�����;���4j��574u��/v���PUW�4	��"��x	�1���U%p�#!6(yf�ǃpq~�SN��Y��ȣ�c ���F��@,�?����ȍ��:i<��	��t	\�"�,9M���wX�f�Ɓ��<&{�/(��j�̦

j�5f�)�ۇh��G;����%��J��3fOWB��*��t�D�T�@�2�<7l܎��j�t�$�1{&��ڒ�7�%�K��B��I*&\h��Jő
����c��	�3���YDbv+	�J%FVB��N(�a�.�����̲'���b/b�=X�r���p�����!�A�d@��1��k�,�PȀέS�^rz�n�<m��5�O=�2}�	i���b��q�6c:&N�,��ۿ4�X�huE��ȋ�������)�����rӵ���������;��?�o��5u|.��B�v��hQ�O?�K���]�w����������3�>��`��s��������[�!���E~�W��t����~#j��Y�Ze��!`q��q��;_@�[��*��;&�s�Y��U��=x�/˰��5����w�ܤq�q������A@�mSx\��'x�7�i�.��͈��R
#0m�I������(*��<��)��FiY���m_�Chǎ\��tW7�����)�3g��D�k���KLr��M]8��5�T�M7��Z&z,�x<:J���l65,a�99s�P�1i:�/�/8WEe�W���~� �S�ǥ�C����\�y�͗��+/���T1醛o�e�jqY<М��n�����c�B0��ʦq������X�����3O���&��=���w �b�֝X��:�޻Q��d�����q��K`����{�m{����E���xl��ɣ��ew���J���K��t����F����\\����F'����\��3�q�N���;?�W\p!F����eB�VŌx<�C[K/z{��8�(�Hz��!Q�v�1#�H����~v�v��zxH*�2A���A�Ji�GIꮀD��8z�ñ=[��k���Rz�" J������b��jkkPR�IS�b�sQW[��Q	��r�?ڋ��v��S�i��ʤY�`�g3�G�����_�v��S�NU����s�pQe�L����H8,fyYDb���G��8�/V�r9��x%c�cO3>ٸ����i��YsQ=j<��b�F�2��F(8�������2I�t*�:vm��=�(�$��S�|΢�����@g��^Ɯ,/Q{j��]�f�������)�$��4�J �� F�N���n\�p]z��?��Ŗmᒯʘ?�L��:�t3&����~�eśDV�T�Mݐ���R� ��Ϗ!�@��z�,�{C\D��{��+�
AuE��|@��nu����ݣŐ�q>c��y��S�!���=^Ub��Q֛.�Ȳ�aHX2�	C�c�`��y=���<	�߻]~x�AU��]p��x�'\$G�����j�D"�-�H �u"R�s�C�qYvz�p{���4���JN��i<I�Ӏ������Xu2�Ξn�r"%e��ciU��0at���) R+��$Lg�:��P/�5�bDukx}!���5+�nNj&Z&d�@�4n'
�E�:ɠ���|3A�1X�v��ft���܈�--7	�)y-v���i6L�p׵��U��{�^c��of+?ِ&\O���i�7UL�I�浘N��ü�%e���C�/ Ln<�Y��yMX�#�F���|��,��0fT=B�^�������#�Σ��[�Hi%2�v�ڇ�NzP�8$gp���1�b��b�6Tc��Fh��(���X�˰/ ,���w��������7��*RP�V�@�T�ǎa��\6�p�O���{ى�:�Y�(����    IDAT���Y�Yj�p��^�&�0&�^��k-qA�#�/�.t���������^t�j,�scҤ1h��R'%t"��#����D��׻�����ӏ��A�W�a��31s���=�O�P7��9���Cq�W��o<�e��c0�A��т�1Ȕc:;\��0yV�2�Ŀv��^a:bL��{��N�'�Q�&�*7%�VQ@>>������c���s`�˱Τ��y�8��&���q:��W�+.��o<x7&O#�\.�g�y���o3��bǽ��F"
���5I��\�B�����Te��I��v�C�PS����\q�$��|��#���?��wi�~���n������k/c�͒Kn�����C�Y�.|]�·�z+��C��/~�-�6㡇��;o��֭���'�섀����)%A�����5� $@ۿ'N��S�}��A� �WV��Z&�1�'aΜ�ߗ�o,���#�}��E2G��´ic�oݏ�Ν+u�|:'.ي���O>'	`vrY���"�oĈzL�:}��رs+b��]��O�v�[�~�}���^���-�� fd���K�K]c3�(�����b��dix}|缺�4�"��]k븜�<%eY�g��?�k`�܌ع.򠺺�dZ���/�?���sѢ7�b�*��ׄ���Hˋ��TS3<͹s��Ysσ���G�?���7��}�M���;n���#U$1��g;������]���������ȏ�߽�b�|�i=ւ���*�}�}kyk�j���8xL1@oO��-�w~�n\}�h[�����X���xkkˮ����ӂ�.]����7z�����X��G_Z��;������2#����btC�?o6.��L������Oa��-�j�Ÿ�����<��ŗ8�Ԅ`I��R��E�(�8b ER�$7u�0�zB���r�A�޴�B)�rd3��%g8/I�I�bR�*��Kc��,��=�q�P��.t�u�(P &ԘI1[#�EYi*+�d�#~�<mο�L�X�^��U��6�߃];�	;��Ձ��#��NGb���ɉ���a<&]v���UY]eE��ww�6{b��h��F��P0�Gf�#Ǣ�v�&;�c�E�Pɬ�����Ŗ�-(1	��R��C���P"��Z�sVL����g�2�n>������v�ri��g�LaBN�NG�"r%�)��g��R����Ħ��R�HT����j.a>�2�4�^�t�G͘���e�58�z�dBA�L��������C�CQ���S ����i��T}�@���(�Γ�7U>?.��"p�e4j��~� iY�E�l�KyPXDs�ba�ǒ�����*D�ڂ�6�^'�2���%�����g�RI�3�������H��f�I�Ɋ1I1ĉLLs�Im*1���N��X�Pe%!H*�l�{x�Ib���=��Gӱf%-��18��k� g�`�#;6|�5TuVp.��y��X�WBg��=,4ϟ.ڄ*ף���a !����<���!�"j��Qo*�v��3yB�2BGh�dt�D�3n͇i���4_�U���t)��%�nw�o%KKl5ո,��0�8���^��m�$���Q�:�Q�����ߣ�;�t�0X���(�K"U��kkQWc�'�S�X<���
"7L�����y�3!�6\F�PK%v<��(��Գ9�Ҋ��A�B����\ԍ7�BAƏGI�gL$��_�)Hb�a�~�k ���VD����W		��$�t���8PUA]m9�K#���/���f&�y�TUk}�z��ծ{��߮��C�t�СC8|���&��)+�%W(B[W7��܍M͈%h>H���G�et�e��Uե�(���-J}F��hk����G�嶹FcF�Ĕ)���Ơ��A��U�<�� rL$�|��d�5�q}4��/iU9Uҏ/�&����*iS[��v���� ߟJ��P@y�'��OV�Dǁ�J��y��:��PH��.���f������]����&���2��/.ģ���:-��74���3f���L
�2�0K�&�LG��&�^V\�y�=H�⨮(���_�[n��U�2�\�z-��o���u���U������_l�/<��G���~��I���G$�SN���s�UW)���/ŦO?÷�.n��6lٲ�?�8v�ޭB�7���q�R.����ēO>���ujx�5�5!�q ʣ&�TQ��$>���Q�8v&i'^[�6}��'hd<1�\Q�����߸��;�Tao1���X��JA�v�9"�	�W|F|>L�Ə�.�00أ���-��Q���@�,�1�F���g��X~<V'��k`��&"�Ѓ����@�z)��Nv�G��6I�!Q����"�������3$\,�q!�Ȣ,R�s[g3���Z�������o��^~�u��Ӥ=�<Er\ȓbу�4ʑ��6���#I���=E����p�MWcTC5\��zء����>���G�6Cgw�܈/��l<��;�K�d�[x��g��Ջ���*��^�l,|�,Z�>��oFt ���r)�5��1q�X<p��pɥ#�.��V|�.��Ѻ}��~�����o��o�K������t��N�ت������U[&��9瞁�7֭ߥ�����V\q��زy��mm���?P��Í�#�b�gb�8�ט`0L��&���z>�D"|��Q|��n���ȻK��+�nBS�z0��RwݕGmU5�%8��K|���p�S����k�6 5 O�!'8��L���GK�JDJ�5��%~̚=	s�9��p�#jQ!�²�����/ɸ�D��a[&
�\c��9��Ĳ�ʿ-+��fdOy͚8Ɍ���#����F_o7��f�z&"�:U
iڇS�2��hɼ͝i,|�c|�n��#���#(wL�;$�-�^�=-��s+�D�A�#�Ews��E��.U�(3J5�+�S�!���%6�[��9�h	�͆�1�}�*_.+ $�E��#��g��+n���bh;�!+�,�kHL�.�L�3�pV�Ւ�$-�J�=�%�uq�P�gt�,z�ɸ!9)He��V0A�u2�����(�Ӹh�:��"���Ua�2��
��uJ��M��j]_ow7b��8*��LAM�C1�s:�����P��Ug&gLv"\�zg�Y��	k�ګ$u�3!��\��Y�i�КV��Dc���}.���z)��E���lZ�AIq@U殞~A�5�3�ii��0��$;c�}�k���=��zU����cI��5J�	���c��I�Kx�BV�H���Lʟe���������Ҟ& ��0�L6a����G!�$]ָaJ�:8	tS���݃��V%��0!`�$ZVD���t1AR�eU���&�am�Xl�]{�9|��Ֆ�'�Ƽ�Lh��pT�5��DƓ��-�0��cѡ�CŒ)�?�F�:�uͼ��������=g`W0n�J�s�P7�fYY�J����&:�c�W�=��O�|&�H��U�S��CF݃DV���n����,#1�vj�����ćןQe��bq�~�� ?��bP�
@UUN>�d%I��=�zL�d���L����V����"(�q���Q��
�Cq����8������7�y�)y0g���(՞���wt��څx��
�}Z�,�#�
�=��Bn�ݿG\�X���PG�$�|�n�!���G��/�;`'z�'��+'������T�x��楀�Õ� /��B�vlX��H�$㲘�΄�ݪ�K=�	����g0��]�������1i�hK*��_\������� mD�H�4u���]�h:pP�T�^1�zV�@_�҈"0�#l�	AMYw�rn��F��b$�����գ�|�稩��w��)�:�k?Z���v�С�
D��w0n�x|��F��3T������7��M�y��`<��SR
x=��O�o�Q��D<��{A�#�	�����`�6����͊{�{^ZZ�{ZW݈Q��~���ؾk?ମd��&Li���W̟����B� �,[�7�y_l?�������*!�z��y���C"9 H;�,��Ք����C0"r�\9�U a����xب�}D:�oM�m
&�N���ğI�k�&���!�5��㜹g��SNA$Bkg6~��>��n$r)�[�
m��h����.��~���)6��������a뗻147�@��r��ޗM"��^>4z#�?Eyy	|�^�z�(2� �2�Ǐ�t�����>��m��K��e���}�+(d2X�x1�y�Y���ᡇ��w�"������o���}m�YϦ��t��U@���յx���q�U�!�,^�:�G??������~��UB��/_����U�wx}�).�1zD5�̜�3N��Q�%8tl�<�:�X�&&M����N=	�/��O<)�|�[��$I�4��aܨi�(����)�$�t��/{���8ؑBA�e�xY��u���q���T�	z��Eˡ={�m9��V!�ӌ���4�I�J�j6%HK"��Cj�Qnt��I�}�t�Y�@?R��M�V,|�%|��G�(-��ֈ�Z�$����=����a��\V�G�#�(��`X_>�2m�ɓP_נ
W����Ac�(̘9(
����T��^�{L`㊠�+��Wl�K7�wЏ`���LQ�''՜�$k
��EZ���09Ȧ��|=�Y	A�xB@��<rE��4ظh��U�%�_US٥BMA�L�k��y� ��>xp���p��� A'��#�$��$7.>$�2�bB��,1�����$s�_a�Il���� ������� E�-�MYMG�	aF܌X9�h�G27^�����Nt��j�3f����5��`ժO�Ŷ���WTWicf�MFB�A(���r[�T����p��i*�F�ԉL�R#�H-gS}grgP��l`P��0�<?�u8f��»��!w^7y���87q��h��(�if�͘|�Lk�1�7]�����K!��um�yH���E��7�t2W:1�9��6URE="�9%6C�
S%�3$&$�2���/�;�~�Wk��::�dJ�S$����"Q[�y�Hp�~lL������[��Ц�ꮁ�0	_��.+�sg'v'ȾO$-��'JڪAQn��eJD%�2�YY>[ӕ�.�;P�J�e�=�� %)=k |L򕔐6d�f�9r�x0�KC���y�WN�OFL�LrXU���}�01v��"�d٩"������D���r"<�%��w"�a`pHssܸ�2Xڵk�B:�V��R[
�Xq��B*_ 	�L�2?�b4��B"���<�`��ys,0GzO&M���Ic��f�{�^��H���4{�Pz9�`'2+.޿}�ʸ(����B*�p���ʽ����0irM��3ɲ�x/-�!K��N(�!N���'F�+�#�.�^�|^x�r����܄M�V#��
�׃�0	�"�q4�`I���6v���p��W�_��&�T����W�ģ��
�xe���:�7A�u��-�J�z{��	\(il�5WL��18�+U�ڪR�}������0r�X���W�VB���M���p�M������e�E����_��G�HU���/GgW�>��֭_��Þ]�q��はݯ���o��g�U ��_��\r��8ag/���{�y�up��	���:�qk�g��g�1M�f&�#�cD�8ttG�j��=|�AJp�0D�^��ķ�s?\x����=�%+>��o��O7�@����R���&�<e�8��=��5��G�9��Y��䰲�B�f� ��ڬ"ϕ�K�>#=���{����������R8cܡy����W��ܿ��q�����K�p���������������]����j�|�t|���@I[��$��/v��p)΢��s=G��tI[��:�Cͭعw���_��t�e���A���.��$V�ی�_}����Sr����o߉\2�%K��S�<�c]�x��o���oSG��eaѲ�ط�]�*��3��NG[3�#a<x�Wq�u�@��'_ŢwW�b����{����[��]%�|���^{���b�xZ\O�8�ϟ���QUN�T`��_����8�ڊY�L�m7]�UUx�Ex�7�:�t���E���N����8r)�@���H�@9)��i������bKɼ?�>%"e��N�^�S�F�Bլ쓹���훱{�:t��C>5�`�!�>U���4x
��`R.�5�e8��S1e�8�݀ƆT���������=����O;Y"����
���HS�Ƃ�U9�ܨ(Ŀ#߀;�HbCQ#��+`)-����Z�+]���cF�Gq��C9m����
1-����(FG<��MX��n|��(�~�C�Ȼ�:�Z��! yT-]a>fr��@w[ۚ��h��A� FY8�X1$՛�vli?���������I�Ԥ籵W1��*��_�ўHg]<s/:OG{ڄK-ʚj7.�G�pe
&�@^���Ǭ��~,��$+h4j0f���z�2��a;���n��v�� Hf>��L����aax	w3�usL:!bĠ�c���{Mu��	�0�����/79ڂF�R=^�7&I��2�r��&��'X�sS�8d����d��x]J�S����<}=��'�<��@P�����N�H�9�@����{����@����:W%ml�� JD\��k��/]��Xdw������ �KBdW��g�^jY�-e\�T��:L<����"x���}�\�}}=rΎ'����K��".��b���A��-`�%�A�d4����f�ډ�̉ȗ��IE.!��=f����?����]�Ф,�;�EEY)�K+��Y�G#�,7k�#�U���o�[3X�hA��|Kd�e0��(XϚ�0�-ǻ�)�卻l�Tp��$ OiV�7S)TW��;)�R����4�y�,E'�I-��4���Ld�@渞y�#��D�;�-GuN!�D�$�� 9F�{�5�C�V� �I0RI¦!X X�h¸����5��sʐ�����Tk�����ˤ���͊N}v�0q�9��At{R�"g���%��"v��H�AI���`q򶊙��Z�m%
��D�-E
�Z{�zFH��7�o�8�[�b��5�w�}$���f�RRaɆ�H@3&i�/�C��t�t�����[1a|#�T* ����P�
��b��12������Վ�^��eyHX|)� ��F:�3��.�MW�CpG��iç���<��?Z'y���;�<m�*Oj�����g֬Y�={����r�(�|�rt��˩��#GԋP��K/�^�����y瞭�Axȋ/�(���Añ���L�$�zT�WB����0y�ɨ����!�\��C�Z��'��Haڬ���7�å�%��7���!,~w^��b�~���@�K����Yg�Euu����v Į����$�G���V��b��Ƈ]� ��r�L�ŵ�~
����o:��|f/�*���q���1C� U�~���W_+N�`�ݽ꾏7	���y�	%ܐkG�b����w��pE6o݅�7lBssJJ+�!q������"e�inH�^sk>�l��\)���^���8�EGK��U��(���>��$��c�ҕH�S�㦛�n�nK���'�}��S���{��������X���l��Ö�F�ABt����?M��ݸ��K$��ۧ^Ţ���z���_:�,�������~�%O����%��_t.�}��4^����CG���g^�K�9������ �1J:-~u��MA(\���>-�6�/8cG�1�G��Q���?7B(�t*M�h�Ɲ-�r!�����F���5OC��n}N�@uI�~ڏ�����z`Z�D��%>ds����;��RR��ÅT�����8ef̜��cF
���ȑ�x�OO`Ϯ]8s�̚1S]a���ZXoCT��6�jV61#;�	ĉŖm{�!A[    IDAT{Z�5��WZR,��P�����aƌ��2���˪1K�T(.F8�G��	�C��EP'7�t��>��6��ݝp�K.�E��3!��t�Aa�`�b}�hm:���f���J��.u-�����ˀ�T��+����I��/;���(�pz�!�WD0�sp�yg"�s���K*(�_�s`m�6���ؐ!;!�[���8Ye�	�9G#�i))�!љ�VV >�{�e���'4�H~ �$�	7ɪ�����A�9�xV�sUQ�����OHF���D��!��~���[���ꑁ �m\m6�A`+�	*�>; Q�&k)~�HيֳZ���!}qʼ*X6�;�2��B��)o>��Omz$�:�g���䢛o*����n Ckf_�m�f'a�;�4�	��ۉ�/�,�O���xj�G��@�z�}�&vS��E_�q����J |�L��N ���<>�0V��d��I�-��Ĕ�����y^�v��V~y��΃]���Y���[�d��1�F� �FB�C2�c�Ȁ�8l�]�s�Ԭ��D�������vA�,�
 ;!�xuR��@�hdg��&觉��r�Tq��d`���(,��PřfvL8�Y�l�<��`%N�$�M�p���T��ϕ�>K��YQ�X�"UV��^74��q�2-v"�K�I!q���08g��*5��Ò��Kd�!�����'�``��B	L@�"���(�|�Hjb"�;\R�R5�*V�x,^:���.;M#��s\��,)��duʲy�;\B"v�-%�AJ��U���t��çkW!��eL�lN���Q�P7ў�$�g�&�"�Gq$�[n�w�q3ƍm@��^z���W�F��DuU�x(t�f'�6�1�~*Rx���,r�Գ�QaJ}O)#�T����Pp^^V)��Ν����Oc��Z���!�1%%���f%����O�?����
8σ�9�G�\ ���;�D��w���3NW5���^I�2�c���B$R��$���ړ��5z��� �.`͆���bь!��R���p�Sp�_��g��L<��@���o��.�_���?
O�š���=]=rt�NEY	�}�-�Mȥ�"�WDH�eW?�L�0ЌHȬ�3�f�ʎ_���~�y����Sa��*���L���,���R)��s��k@H#�^_?�Z;����\r)�:�Zp���Sg����8���Sغu�<Q|�AL�6���fD���+?X�����W��c�y��6a��*WkOm،��Y��.\r�����KQUQ)�h�H��q��s0z�8���؏��}	���-�߈��u32���\��^U	���ނ��{��xi�*|��6nBgW�~��q:;�XU���U\}��ړ~��+x��[/�7��񃿯����.����V���s挺��k1atJ'H���-�����hiu5ʫø��+p�������p�[h�DI�Z���O?]x6F7V����O�1��n��^��>�]�ўV�ہM{ۑ����B"�EO7mʍ��8l,�E(,Bq���H�!/�(}m����؞�qx�f���+�=ۛy%��D�je�MP�ȁ�
?N�}2�9{G֠��(֮Z��.��ڬ30��^����,-7Z:���6K���ڜܘ�i�?AxV��8��P��ߧV:c9����ǅ��ᔓO���p��:%�!�R��Qm�\
�2�t9�z�a������(.����:	���h�	�A9!Y��k���]��~p�T>V��yn0��@�}��l=o�$�7尡VŖPu
l]��OY��7��;��[	A��<[|Y#�)�/{�7�&6����;��s��{#4�G�$�#[�捖�S�L-���Ҩ`Z�F	��7Ҽ�a���j%'�`	C�rI�A���lC<L���ʀD�T%��M%VU�\vmR �s1�t��Tj'a�SpCf�$7RS6mb�i�eAC�b��hV�p �z�|�ÄD���t���$�Oȃ�D���cd��� ����v��x��N��4|����'�v
�fu���xB��2��"dƳBj@&W1jR�8]Z��AH�]�
���g�#��H�r>����e�;=3�[�cs�q�W�=ޕ�B��dW%1�"���x�����؟�@���9p�q#e0#l��%��Z�ɔ�1�U��Jؐ8N�
'HSrZ��K��Y0^�}=^���-�#��T�i�F�����P�0�,uJ�]��3�����T����s���I���[҄�r�c`:v`�HȜ�( ��H�OPVQ���"���	��5��p6-����]�-�Ǚ���o��y�r%I�M'��s�ǍT#��R�a"7�繝��p���g�C�Qc�$x�e��@T�o�����<�d_�~�b�#�g��5��\�)�`|r(���Zōl�\�A�[����e@t*HY"�&���$̲��Ɠ ��V��*�����߂������sϾ�����E8v��n���#\Z&!����_�KF.K2���t��&�����ea�Ո����&NИdg�����]��k?�r:9[6���J���bu��{��!l`#욒+AO�tR�Bp��a�������'M���T��~�m���B9�$r<9W�l1,v�X�`�j�F8`�U���+���/v����XVh�ljH*V��N�׾~�y��(�%���ko��g^\�#�]p����66�=eŜd�]۷����"�������lZ��@q@�%)���d���p������tT� �$�'����Q��~�r��y�ǃ��rA���%��X��'̞1K�)&Rq�m��O��Mx���úui����٧�?�1F����Wb�ʵ�b���~̙s:�>k���z�PWF^U����I�Y����/��矍�.�X�����0��{������Nbْ�r�w���|���X��*,Z�G;:p�M7�[wކ��$^\�Vmځ�:�14�?%�	uv���>@��� �7O������%2�-�7�����ǟX����Rq�P(�ޯ^�b�ǿ��ƫn��"��ك [����U�b���Q;j܁ ����r��t.{���e���/!��ǌi�p�50���dT���^�n�R��:�:X�ҵ_�-p��7\�h4-<&'�H-�b�� ��TJ!&���~����(��c��vx;z[�r1A�E�G�ȶ�P�p���Kr��'�k�ĕ.���碐O`Ųw�y�:D���6e
�*��g���bi�rq�2��;w�@wgH�>��99rj�qwL$Y�ۃ���c�޽���!�֍��/��s�'i,�@<E�Ј��$a��l���4�9/\�J|���.ބ%+��f��;��#��"�l�$,� ���Zސ_�:�VPj�����:t��6�p��ѵ��v�_�!L權����ϤK/K!��`N�\�#a�v�\�}Ʌp�=h�iG"K��S8S��+�I�"����p�تX�At���0XWࡊ#����ɖ|�00b���B\��KN���xצ�=@�UwvZ�A�� �L�o$F-�H�v�Df,V`W%k���3a�p�i�&�� 2'��5��Ov�e�	�)&#3&���G�d����|�����	T�.�@�ץ붓A��K
�����'�-�$)��2βǃw4�z��9���l�G�Й`�[�[����a3�B���_'�v���A=;�L�>��Y1�a>JY=�|�ENg�?0�#����]���Y�!���4�W�`��Zɑu}
���"m>��Ngg��W��� J��^�
�P5����,*�e�f��N�:M�s4!�!��ɨ���l���*I���[�)����/U�������YU�5&�ڙ�yRb9���rӵ0P-�e�G���5����dë ���Q�,_D�ܴ`t������j��d���\�)8�P��&,�;�����	�gJ�	IV�",&����mu0�{?m�Td�>����:s�)";Z��G�LA������ʿ(Z�w�8�'�l���<+Q0]�deX���g�<��*!�)���(�._���Di��e��R�!)s������_,H2���K����+p��b��FdS�3��/�g?�w��F�BUu=Ǝ��ѣ?ٶu��e�>s�R��.�$��~P=���Ғƍ�SO��g����:��ءommǚ�?��M[��b�+3w4�ƳsVP܁/&���u��@ǿ��UJ'1y���G1k�LU���I6&�xێ/M���ֹ��(u��}ɝSJӖ�KW��/�Ͼ؆�(�C)%9	��0��)x�{p�ٳ������;�W��g_zM�:��^� q�k@e�8�������!�!G!�X���|r��2�$���Z��1ޤ��_b���	c�y�,p
fSU����!x��.���{�����Ҷ�V��Ӧ��t��g�_~�̘rRTet� I��.����;����	,}�}A�2�N9}6~����x}�2��b���`�|�#Rt#��O��\��S&a0��ҕ���3ω�v��W���/FYe6o;��_x�>X���|���ŗ�G�@G[+�9(�����!z�{+�x�2t���[oƽ7݈x"������ԓ@�`B|�x�R9�{{0��_�������e�^����Gc��/ϝ{��W���(!x�Ppny�/׾�h飳��������z�;�n�Z�߰{��g ����*u���.Ăy������K���O�3�V6hp��z҄�j͜<i�HKNBC2l�S�# �R����?ޏ�[!㮄�_%�5jlJn���.��'A�6�#���绰m�G9�(�d��v���Ļ����Q��U��>~��3�1�ÙÅ���7,�)3&���0�ڇM?�`o/&������͛������knV@2}�L\��*444�[�@�
l8r��i�D_�]{vKW��s���-<:��nC��{Œv#n]q։��I��|�.<��CtF#�j��t�ÏAU�(���8�)$A�o�Q�a���ٽ�--@gK�"���߀��l�+\���J�2���L%;oȡ�� w#�ץБN� θ�<̻�8�>4��1M�m��0�ª̶���Ą�N�3�)���V:�ɉZ	A&o��(Y�4�G�9�b#�'�B�	 $	?�ު����H&d��`ᘭ���Y�[�^�&)0R}�9��|1����K%��*����{�x��_�'�����f'!�
N�d{��U��`�-�ϗ@V�U>�"I�$T��>�w� ��^���e�,�K���X�u
�qq�c�$�<X���0ؐ!�,lWD�.	�!湛���!W�	���I��2�e���wB��� SI�U9f�Ī�%�E�Έ��id������'�3�P0�	�`�aTvg�Eb-�Z�T֭`�F9�V�q&6���0+��us����*7j��K"Ad�q)K��������@���)(�:lLtoe^��7<o�����uK��m%h�9X�9!�g��Ύ�p�k��1�{�J/ԏ�h�ˀ��<3�������7HS�ά��9iا�a�3�%�e�=�8��x�����M�p�x��!�؈I�ԍcBo�qΐ;�s�����N\��n'9&94	q�Q6�D<,��4WTR��3���|��q^�M2`慕�Y�>?��X&c;L##i9�G,C�&��4FV�!�Պ���E��K�>;�<&��>��L�,��[@9R�D
i�{��W���܊��G)qa�C��|C�	DJ+��8��v:�L��CG��sۗJx/�eOg��Z).��NsT��¸1�0u��;�LL?�ͭ2Iܼu֬Y����LJp+���s����}U��4�x�}�I+�n=7�"a��:���������^z)J譄�DU�}@�ev�8cq�&�k�s|ѫ��gJ���0r2Y��؇�"��D4�4y&�Q��Y�o?���?S�b�O��o��^X��d{IӠ��l
�rea��{vlCs�a�3�&�Q_[����2v�1Y}c=�����pW���/<w;9�c�ߟ(�¢D]�%�;L�\י����AΧ[�!��}{����&�|���� c��A��z�T�,-�����g�[�Qq��g�z~�دQYW�W��7�Z��M=��R����>w�X/�M����
.��D�9����x�O(����;q��#
b�������JF?�Yg�����Ξ���QP��4T���^,^��Z�݃Q�u���-׉���K����q�s�l��T����&���?p7�/8C�4�%,{M�����y�����_���C��Pp-}��^}k�ϋ�K���R��C���V��>|����Z����#R�5W����3s��O~o��&J�G������?g�~
ʋ�H�p�p��y�(r��I� ��i3>�l?z�~�]%2����b�3��Y�u�ȼ(��XЇ�{�z� �C=h(���@���hۿ�v��#��IS-<� ʫ�QY]��d�=-�2u���J\0o��BȤ�ر}+�|�R��$��7F$,�����ۋ�h=��b�_|�8��yzB"�y�>_<g¤����@�5�}ͭ-8��&���)S$�G�K.dL|X����G��xb97�I��WW`���(G�b�D����.=h~���~�A7�˃�o�����AwS����[�D4\�ʍ\��M�s|g5����j�+
4��ˮ �;i�S8\�9��s/�G�G;[�!0Ҕ�?3%���w-c'�2l�;VdH7��Y�$Z����GU��@�	O.�\:i*w��h
�m�3�٪V�ؘ���
���b �[�S\V����O�Y�'��$;'�O �m����W^��dd8� �$�m%kZ���@Ql��`��Z��P�Z��dL�ѷ�"�ֿ�	3��snv�۪�RԒI5����u�J�,��O#=UǏs(�����@�Qѝ�=X��%3ʾ��x�FɈ�s\1ˆ)�����Cb`��rL2P��dp��ň	`JQ��~��$ikY�2;A�q���j�)W�b��*�q/[����o�Dy�:K㜉`4�/x��	0�ټ:_|�fC���V����չ��@�(�ء�� ������r��b��z�jl��L��/��(Q�������q��kw�l�Lb,�LV�� \�Ҫ����{�Z����tP&wv7�x�݆&�5��cun�����9q��SR�cဢ�s�����Es.�5�/���c����@�$�C�a��'�l�	�����4H�L+��)��Sǜc�w�}]p�R][�TV����v%7E��j7�z��� >k�Ӆ|&��H0	:8�rÕ����1��V���y����2.,-�Ĕ)�p��9��I���,RkL2���R��0��$���K��(��`d}��rN=e&�i��ի�*L/?SP;¸D�6�JRF o}�C��oH��+�궁���Ĺ�N&�����Ž�~ӦMG6S��e���W_ő�G)��=�b�y���!��K#U�ǌ�Ƒ��>ڰyg�M�n�t'�C���igL�7�s�%�U��>�sU�4�3ӣI�	�"
HH"��%�1������8���Y���`���L0IB	( ��2J�0�<��9V����{W���|��^KK�QwW���o��}��������VVQ��9ɭ��>����15��*e��c�voO?�=�\Q����2%���ߛ�ԜڷÇ_A�V�����d(��Ţڙ��ׇ�C&�/��^{����&V���N@L
�A!��x��{�Y!���7nx�u��2v��r �/U�}���Ï>	���i���\���������wމo�r;���~�y(/��Z���2�O����+����܎��/���!x���!��O{߸�6���`meU���+/�{���w���DK˫������;�م4>�[�'>t#j��v���݇�s�u�U�`��f���w��g>�	\z�k�R��k߾w�}o�P�?���.����Ͽ|�T0    IDAT����O�!���;���G������V�?��ɮK33Z�,�C�8�tu�B~d�|��p��<����ރ��4�	�Shwlx o��2\q�E�E�d�L��n�g��t���E���A,��hz�h��5%�-*N%l_h��g��a-��r1+���R����1w�9 ���c#�=��!��C�� B�(�V0>1�7\�:\~��8crL6��f�=�N�:�ՕeE���Jf�L���Ռx�t,x�ފ����aju��i�ڔ�i-鞴�1A #�}��C���$�#_�}��P������t�>|w����-���#>8.G��h���|�AU!/�� �1
����
t|(-dqꥃh.NM����t�ڵXkSD��i
E3T1�2�:�t��&`'��'e�t*��/�DNC���֖Q���L���I�� 0@Ͽ���H��`q�s�o6<��ak��1��[$7��>�kjUG�N�(�&:bt��:mjrT1���R�F`CA Q�-|�,X�4�FB� ���>ǭ��6<�!p߳�sꀷ6��~�kd����v���4DX��(���<��1��l(�~��g��Љ��c�bBZ��n
j(0暻߳^��z�7 �!�"݆�f8��Vd�bvTV���R%��*`�Es膺�,6A���h;�ZSn#���3�Ü�0fQ(HL� c*���N<Lrm�L.L�{h�LJ��1)E�B��V@��4��*����l�s|fy�ҝ��6-��m3���b�JA��{����+�MC��u���e'����d%t�p'U�il]�_��m,��	��!pC�u��Wwo |�B���W���Y�,����V��E��,�Pǲ��HJ����a�0q��Y0ʹ�.��E��CpM�i|��6D}���2����oK��dsP,�LD�.�m]�e^�k��n�FX��n�=ϫ㲍���u����3j�Jbx��(�u\��Jp]q V/�طu�O�/����UD�0Բ׏�ỲǤ9s�ƽ����J�$�!|���>p��*ܬ���_��5|��_�����I��{6�Ln��6���S����T�a1�p(%53W�z&�=�z_�X�\q9vLnE�g��EfI3�*�g�����K�J�z
��X;wO���s�R�١��+��m�u�^�w��@'���O��_F�TB<�Y����L�ߋ���Ӏ��g``���<p���?y�z�;�2�<.��|��g睵"Z��&����N�z�qrfI.C�P�ZK�������s�٧��8�p�k��pЋ��Q� �]�2�0I�&g�����k�K�.Rij����w�ܭ���?u�l�H*��$�߿?��~��������k�p�t,��&
�y��x�l���?������D�������x��s���������gC��ՀV�ٳ����p�����[�����5�|���uo��H?�����w�P��&�����nx�����n���~'ݶX�1��ޟ�����}��'>�i\�v���w��K'f�"2�k�c�Xۋb:��/�����q��c!Sė�z+�}���Jz���.��O��������=|8��y�?����	F{����`��F�OnF_��ǁ� �cd�_p�>/y�a���K�����	�����׽o{�5��A�L8�)V��8|� �M��'����c�BY9�O$��%5�.a�Sze�H�5W�!�c|d��*fOB�S����©�(M�S�jZe$B���6�#��"�ka۶1\x�Y8�Ha��14U�i�>r���߇�Qd2e�޻�x�;p��stඨ��Q�|׀?�J�����Y<@|Y���jF��;&e�ǃ%�c�^m�ӎ�\�u�cx��X��P�&��7�D��<).��%�ۢ�O h��@�EB��A�������C�Ν��Y�ذ���Nn��6N�ޚI/��=�m1a��)*�tJ�{S��Ej"I,dVQiVe��Ô>�r[��4+ޥ�k��a^�?*�jdh?֎���e����)�J�}-V䤲��/�`�@r�m�����q��gu� {s��}�������4*�'��l�u�'�'��N��Y��7_0� ;u����D������Ы?YN��������\�|^��\��u!j�sŻ@w�XZ������66@�]7D�Xskp�8�x�6@�D�g���4�/����o�#o�R00>�%�m�ᶺ��\&���*�
BkE��_z�9I�����L�bd ���d)c!���z�����4gY5��	y�����g�i��yQ
I�cG*Č	����l]#��2��HK�ͭצ�6e����'�lB���k@��p����	0�8�v�x�b6![zl2��Y�\�ހY��EO>\�Ca1�3��u+n]u��͈\��z�u���1i���*чl�s>�P���Hw4T<�����uǤ�M��}����|+σ�˼��84�.�a���8��Mۆ�5�Q�2k��|��z�b��~FRQ�f%*�峈���a��Fq��C�6�t`#��QA>��T2��|����{�0�
m����O
/���ر�L�ر���� �����e:�6_����B
G
)����,�RD�#�i6�\Kl���ׇ������3��Y�j�����hMm���
YKBKhM�{35u�|F�T:%Q�� �h�����
�T_J����aQ�(��T}ppmo�]�܃�Ba-�()
��,.yݹ��?�,�ٳ�=��6����㶻���rQ���T�bzz�H\.C�x�<��Ve���q��UGuX��}��pl=���0~�k��}�R@�*iXb���Ie��Ф�"
�٤-��
!��y˖͸��{t�>���㒋.D<F�\F"�� [�5e�/���ȳW�W�ޑu�_�����^�B1�'�z
�P{��Ț��Lz��&�\y�e�u�>��fq�w�{�}_�C������>�쉗����˘_��^v�m�r�99����o��F���hc5�QB�?{S���w������������㕩9�8 ��]�����Û��fl�9��l_��]��?/�.����7��O����=�ݣ���?!x��ӽ��;�����?����b�~��m�ţx݅���wD��#/��󷨖JZy�X�����AŒ�6�)N�/:w?�|�58c�fM"��&��B0�?�Z	���)<v`��(���fn�&n�p�t�yR
|��N�f�f�C��:>*q��F���h����i��!�e�B�Wm�(���(z�\ULn��=�14؃�?G�Z�@J\�c��ŗ�ñ�1=u
�l������9$5᳼W�P�P��P���,pR�M��h�P����S8����%��{���o��ڹs��%���g���|;��􏟅B;�N0�6'9�6�3�i'�|���|55D�C,�*��W�p�$�s'�&7}��FRv�]����i
���m��{e=�¢L�k4zU������W��^s%=q#*��z�>z������ɈS��\�g�5�:N��с�\��qf�EA�?:�4n��b&���ą���U���,[�����(w�?Q���y�2��\��ޛ���u�Y�
d��\s�bd�ּ����n�\w��U�,bAC4r�m!�ɰ���"�z�������[��|v���FUb���Z��~��Y�[q��C�����Q>֛�.EҺ���v�Š���Ϫ.�����Sa7-������J"�3��;�!E�|}+,4�cu]�J6���kݮ&;�2�
�6��r��&C4�p���R^��!xS,�"��=�O.JJ��@�h�Yz��J��O:
�B��SnuΪ�W"�S�;�AW=�ƈ����s+�y�[TvcA뮗�k�:r��M�M!l�u\ӹ�9�^맭�a��7���w�4�*ǵ�A�)�r�jNC��k�=�K�8�#S�.4%� �'6�����knE�v�r���lZ��5>f/s���{0����p��ה�/��FP��QZ����4	���}X>}\A��E��E�T���X�2��W,���Т�r� �F)����>���}7]�͛D��s���}_�ڷ�$(��������&�.8�8zz{O�Pm6�+��{ﴥ��O�y�vP�eՐqP�g4�wt��{�037���R�	�iiF�eSvύEe���s"CM��J/QgA�|��$���:�{�z��4�H���	��)�Tg������z�ʱSx��d}�YZB�ZVH\�^�ŗ��?���b���4�BX]]�wo�7�q'�Wr�S�@�Z���S�9�h���{�����"2�j�:ф"�V��B��:������	ˍ���*-N�}�?9�O"���*�=A��j��� <�<��8�7��شiX��U��}.���wʹ1�/c%��/~��
_kyȕX����މ����`d4���U�/.��&���HH_2���Ѣ�e�́���?���y^L��|�{p�uoC4�Ľ�>���_��|^Oo�lQo�\q��g;&{Mh�j?�1�w�8q|
�{�M��܄�x��Cx��#X�N)�m��Zj�.���vn�a���Ï�~<�Hin��׿��?�������>����!��������O�y��O�l��5g��AO4��y5��bz���o_@v����^�� ,�+�2r������d�K<C_�gl�*��Bk�|C�PA��	̧�x��x��
r��/ʥ�
3:�p � )D��چ�UJ�ZC��I��Ϥ1}���E�=U�y���P�-��2��*�0xz}O0�R�V,�P����>��]{�U��ګ16Sg���n#�_��O?��o����7�x��GWo�)�kMDC~��P�mX�ZXn�bK0�sϿ����Q-�Ъ6������4W��w���K.��{Q* _��;���%�Fv"20�J'�"���<"�|PPʩZ�����H* O��B�Sm�!��d�|�˳�4�d���3�Ąd��ɔ��1N?`��W�a��<�EoaA����Z���I����������9�u���M¸<��8����eU�`"�6��In�W)�s�U&vC}L�RZ����2��F���F��nD�Jb%�m��F���,2���[<��y�4�4y�<�c�:=I��|�F�h���ˋi2�tԐ�L��r�v�f���9�FBԏn7��m��"�rI]����&�N��S���&���fZr�qT�Td�P�~gժ�M���e�?�~�Ud�!0�װ8פ�;�!;E�M�l.-w���Y�v�o��˙�7��+>X�7uDER�I�愐u�z���]�5�H�6�7�q�p�K�u\�H�]�Hb��i|�ke]�4��-![������� F��DZ�P8�
y6��p��s2����� 6 ̬q�
p0` kg���E%��rt^��w��n�`�{�Ap?ǽNZ5u����_����-2���g�k�G-���P"��t�(��̾blo�3V��Y��o� [�06�������6\hX�`wH���zm�����;:�k���t{����5 �Y��)}���ϳ!0�;�m5>a�C^��N��Cem>".,��,�7�C�(�KjՂ�A{��O�&n�����/��?�_���ar�C(W]��⠾��e!����'��NQ3ғx��*:�:"L������F
F�����.8_�Z<������XI�ɉ�띃&5��y}H����3j;f����D�kA�|.�s@�Ki�����׊߇D*��Q���ӊc�@Q��e�波fQ���(e��4p�E���ػ�}ޘ?���,n��v|�������꬚�Yz�062�}�iL�:�F�"�����X�J�J�����^GKS�7:@qߡ�
Q6o�y��b�� Ɗ��1���k����1U����G=��Z�4O�w��{oz���<���<}�y<��a�I������Op͵�G_?�.���F����{<�6*�2>��� |�1!}�)���?��{+���a|�[��J��f'��7��bc�Q���w�C��$�����?���{/�+�x����>�A�1ڧ�U�mH�]k���ͬbhp���>���s��S���������ţO��]�������^��i�{����}�{y�S/~�g�d4�A����ҋv�w\�M����)|��^9p��z��Mo��PB�:�+�U��a�%(�8}|�J�^����0*0��Xb=X̚��c��7z�����x�I��hW�Y��p��h2E���J>�|@����shU��k�-����Eu�@�N�y;(��G��O�>���Ɠ�Gp��a�]���t �<<:�P�w�Źe	��d�O�]��j�H ��<��P%�ڤ0%-T`ye�A!����<� �W������EL�TB�E�����mx��Ch��݁���&���r7ufX6���[B:!
��#��js��z�4:�Ex�LϬ�!`:��h����yaaUC"�lt.�I�^;R�R��h����o�������:89Z����:z��\y����Mw��+
�c��V���Yί��7p�:��h ��'=��~��G�)	r�qV���Q
h�j~v�����'g�aj*�.��)�{�uY/T�f�����rAFn�t*��l mC���U�ʐ�T#��\��/�_���ES���5@,�MQ΂�_]��� ����J�r�����t���A,������4��H��j��q��˭O�I] ���LS;`P!��� �i�,I[Ʒ��!򾽖�a0z��BD:���0��t`�fZk�,�DTp0��כ��Y�r,�b"(�(�b�M���\?\��$�5i8::���>5A�N�&$>t�i��TQLlhtj�"äYg���=C��Zfm<����W����)}������j�,��BN�:U���V�4D�
�m����C��d�
;�߈���f�͎C�������#u�\zVt�4`�=�f�Ar�(���}[�k�u���Ʈ_!�a5��n&�K���/ol��>�(]�yx����j���L��`_�|>�lQ�`�5$��А��h	�F��*�<��(�R����̰@�F��F�TQ�ٮ��F=��ާ~7���1>ү�f�ߐ�Pn1m�؁�Va�c�`7͐��zx�O��#X���&*x�҉�\&ԩdZ5���1�B����|v��-[ә�y�ZD�:�H �T١�耆�G���+v���b�I�WS��}�ӑ8�5�&��2�@?�F=@,��k uA�3asʡA��G0чP���W����i�5�9朻�����ۃ@��<X^���������:>��DRMN.�E$�UW��#�x��p��!�+Q`d�_|Z��у��#���g�J�6��!�A�K�]Q�;^c�+�I�JH#S3ժ��J����	�&�s��n!�5_9_G4�<���Iϕ��G�h! ��B� T*��ګ���W��R���� �k�af,��ԓ<�����Ï����h+H೟��}�;���⎟<�\�O0�H�G{&��jagl���S��׀/��o�+~���Q)0:2��~�ݸ�u�a�?
�,�"�����ͤ�����K���'�E6����Jem����᭿�����_����_�2�����������Ƃ��N�#�2F��\p�&��Cx���{Ŏ������#�>��BsP#=F&����O�	i �7�3$�o��|L7m�#?o(�\͇�:�G_��Z9�b+�[-�������5�&��_4[�����1K�9�����9dW�P�̢�_C=����QTWf�JѴr�@1I��?(nn,҂br%_��;�k���#� �'Fq�Gk�    IDATÂ�<�����DLLL`߾=*���qॗ1���b��VֲBX��
er=x�A����lx��ʞ������m�Ė�{���P����A���	S��A���LQ
�{��Jn�@�'�0���%�8r3�@n	�F�4^n���s�fSpol�ͣk�ĂN���:m��<@jhH��W]�FЃ�K���+U��vиKFeC�����Fʅ��-�_(�)�D�V���t�&��"���p$(��]nR�
�@���*'`L'eA�l�\���Dt�Ri�V(��B���x@�~dy]j�}��d�фL�b��~����n�)��7S��k�m�Ҧ�Y�c�kp6Ѵ�c�J1�q���QR�,��D�B<��i	���6�݅.M�6ۖɼ+^��JW�V��i�/���`4�;Hf=p�٩�j����;�E�i�u��˦���fUM��N�b((|�*����;[G�(+��EE���k�_<����L"�4jR�x+|�7�k��g��ŨiN�]Z������]a��]����r!�V+ISD=Lќ,E~87]6>|�������+�?�~شf52v����bUG�q���u�Nos��]Q�͵pz~f�����b�6J��H�[�눁��p(�-�F�5,��ߎ���T�
)sRss=J`֊A��IC���y�v/�M���X���3��b�hKa�b�*�?���?�>�iZ�G��V����>g�L�Gm`& Q�]
x��F�^��E��t���j��;��VUUY?�!����U!��w����R_Լ�zHѲ�Z�&m�gUЪ��{��O~7���<1"�r��G~_��o���i�t��)�@h"�J��(?dԬ%��%D�45��&�|_��) e�z�����g��3/��
3|��'�	<���`1	F�3�����ب�z3ף�`<j��:BX6���.V�Ѿ���5K��̸�� � ��U��B	�R���� �YFqaθ����}x�U����w��D�^������wo�M.CWy�k��C�\E�'�+_9FF���O��WЬUT�0�Iz�:���+Y��Z��i��7o�~�5��o]�I46a���ڭ[��Z��JSZ��^3+E�B����~x��jU�NKUm]�r�Z#������
�
P��	��K/�5W�۷�B4��z,~E#!�,,��_�/�=��Ss�z��@8����o��R!?y�!<9�v�� �MT�����r�fW^y�y�[��������/E��&���x-�;g?Fb)�ǒ��IY�4td_#�ZË��Y<��A<~�=�4z��Xo��z��~�g���O?���<��������_��^_�w!O�H}�6�l��uo9��;�\�>�<|�0�9�N�P�@! �VK�ey ����5L����g����;��d*b��C���`�?��7���r?}�(�4�	0b�|��oZ��ׄO���@�?��(���]Ά�ը��,��^TXY#����q�LCym(f�d����ޝ0��N����I)�2ݱ$�Ѷ��ؼIH��v�Ã�D"!M	�F�q��N��b5�CG��1^"A��
Ut�1E��b~yU���Ilڼ��aK-�[~�R#(�(4=���Hģ��˨R#a�kv�lhB� r�,��*�����bX�^�̋S(-.��2+�����j�7�&�<@����\%�4n�F�&��P7��.8:�}��2t��/E'�����ͺ4F��.T4���kr��Í7M��&/mӋ�2�"���9���7�욒�Ñ�x�##C��P(���Q,5.M<p����A4���˴,5
�7C2��e�ҘA��V����'�vl�ύ�5�~�#��<reo��d�g&��E���w�w�SǫI3�k��1i�(Y��)�T�u�a����uC�( �OU�f�ɯ�m����6㦙�s1��,��l
.g�h���b1�(=J�����r���J�N����=6��6�>sC�FS��QCc���.�Ѫ�H�k��%S7E�-bI :�b��_��v��m��'����h*�(����X䄔�~�x��3���b�;�~�c}�Ɂ&rf�s_�Lνe��
A����h	g!%��&��An��Զx�)p��_�ø�lG92������FKϫkY�Y�4l�r\q��w2�5
n��m�]�WNVG�YoƝ�)_��V��ܾ��m��XMg��(Xm�gQ����Ѯ�>��Ym�}�.@bm!}�n�k�&��#5�r�2{�9f�����V�>'���1H�	'4��z��&�r����m�GBr�/��Op�4b���Qwd+��\i�&I�{ =��B���w��vLNn�n�hi��?�$��Ew"i�f.��v�|߲��L�_�#d�L�-/�
O![�_�h�L�LZH;�k��+۳y��M��@�Z�����������{ H��x���y�tl���Ů]�q��-z�ڝ�
h�8�dB���鼳ϥ�p�"WP��~�HI�KyRg8H
�� ��aM�i�m4�9$ca���}��{IIެ�:�a-��-�߁o|���_&��Ui�1��K044�G{�|Y�T"�@o��n�r�r�[����H����4{������;��Ќ�0G�Yr{��HR����=��9(*��H�$�z�}�BZoD$�ggt}z�G������sExAt*E��>Lnٌ��!C'�h&�:� ��2f��Ih�(��A��$vm۬=ujv9%��h�8@�ˢ7ʡN��z�l�=g�C$�ZzǏ��Jf�v��}�FԹ��2b� �z�������H*u/��<w���VPny���ͷ��'���W�[���3�6�]�4�7߸��x�����1�/���B2B*�ǖ�8��p7>|��HR~���]�+���i�ԩS��3Ocnn���G<փs�:W\z%zS��8�6n����a�<���q���P� �ބ�$�(`ż�B6�"g�*Dڈ�M1�E�ŦC�UC��A*B~m	�Diu�R�)t�V�vh����4��GSa!
mȵ� KS9�lKh�4&bR@ٓ�G*��M5��d4T
��� ��1���B���o���!���i�Q.���oɞA��[|a��w6F�7+�P����P_ z�2-7gB�L��I�!�D��� ]�(��!����CS(�̡����QF�C����i:���<�;���ʟ3jG���+ca�/�9�I*�Ӄ�/��}���r*ԫ����Ħu��֮QG���"�c1%`j����fo���'���/�A8A1�E�UE<D<���q��1	����9,�dp���V�G���?)�G��Zc�C�<@$���� ���.t�k~z~�B�z�kjltYǺ릹�O�m��f��9�S�r�iSYCS6�~U�4\e>|om�r!N�B�E�4CI�����p�r��|&tG���D�\4u�ڲ�[�eP�4���x�� q!Z�ڤ��S'ֺ�����4=�bh�}J%%�O���$J:����h8��I��
+R|A�y��x �}Gc��C�M4Tp`܃����k��i�7>U�=�\�c�H+"�����F@Ȁְ���3'������H�,�t�l�)5Jzn��I����Z�뿮@'RX�G#1�r�����Mp�hB�0���}�FC�[R��Y/r��x�l6&�¶�ʽ_�4�����UMQEPf��S�e�b�V�� n|M6�>Ni-�,2;�VB����{�"�a%���<���0��`������1M���-��1��#W:e:tfP��Akok'�ZK|ߴ+���4�ؖ���&I�\k�
����!�aG&�ۆ�Y�aC�j��1ٕ4�Z>k\���i�b���� O���3�qꐠB��8�٠�4���ƦgB:"L�Nv���ВZ�&�.PMȔ��5�xZ�Ƶ޳���䱩7��X8~��u�����O6�ȏ̢4\'�#��m�������KNC���*�q�U�"(���CT�����T��E�Ը4%&כ!�b
X�z_o�z	~��V��+�3c _@._�iG�	�,,�?�=�4D&����>I�K��'�)�J��qx2Ʈ[p�%����ئ��q݉VR���˦�Ke��ƺ��X,+l��%]�:�ᠦ�J��Z�?CDC�sh�a�Ո[r����l� iE/���W���-��ͷ}���t�~i��
E�k�p�����g8q�X�Ac�a"�}�:�l!#�h���4E���xM\�+C�!���y(V�{ɺV��.p]+(РTל�GtMLsGףx(,-���f�P���76�P4�ӳ+(�k@�Lv�<��j��U,{�S�ϡ?�j�)�y"\�q��=��6��2����Ec�V�?֣�s�H����^Z�?��Ƞ��XO��%�baL�8�p K��j�X�p0�(3@3���A��F�Vњ���4�i�ҳϾ�͗~����{���i�x�-��������ٷ��6#��:���|������ކ�&R��pr����"ۨ*2�B٥Ez��P�U��oۊ;v!��1���@�@�Q��!8���e:�{S�xC�	�`����]�)�'�z�^�!Q��&`g�1�͡����8y���C�UC��D-����,*S�w8�(i�c1χ3���4՛�S 7RN�+�`.S�;����0`�A8Ef�C��� Z��9R(:^��!N���^�#K"K"I �7�J�p��D�@�RC�����i�| X���ll>���Q��r3y�m��(�!,X^�"}rk'N��[��Y�h�4��5+N]��s<I���2BbM�Xh8<�d�$ܹ)u|�z�p��W�+.C�,e�Pcp��� �4_�Ym5"<$�*���CJ&b�u��d�OF�xQ���Y�ͽZ� I �c`K�*ӟ�8c�VLn�@__BM��J��W�M���Yx=!m��|^vzlz#�$�
L���b�X/&'6iBQ*�������
�VP�(:����v�-��G���f�ˆ!Dn?Q�F�H=�q�%�m��<>3�$xPV�p�fخ#�c&�>�N�z���jG�lG�*m�k����_�X��(r����=ɔ^[HM�%+@o��g�"���Ȝ%���c��܇���:�O��y�T���+(3s��D �3Y�5�(���e&�L�#��m�h ��9Y�sa�>LC@{A��H�
��d����X7�VIlg\�7wM��M��Ն
�F�]�C�|���L�b�A����J�c�Di��'q,�L������'���n<��3Ң�	�)μ>�}�׌�k �T�FS	��D�Zcjz�[d���r�C��?f6'"fѪi��K��)�XT��&zl�����z������7�M��ll�F��>6nS7&lBh
R'�7���2�v����ma��jz�:��c�,� ��,�Ig5�~;�����%r,=�-�y(e# t0H�Ѡք� q��	�I6����R;��iK-P�j(c,��ZV����]H��	>�A���UGd(q.qYT'��@�O�c���2�F�ql��҉#���[Q�d
�9�P=�Wr}�R����ڪ��ˈ%B��} z�H�Q)���R�:G85�vݘ�qHc㧉�"�Ex�Z� ���Q��G�-f@,d�/f�z���CS�k��n��.|���ıc���\ ��#at��>�u��������s��#y�=�Ll���w6�B�8��}�TzN�Zs�В۳�c����a��`E���d�0���E��Brpb>���P8��ͷ܆�o�3+i!�jv�MsY����k�<�aiyA�/���e������b���_,]��Br�q���4ו�㬀��a�!�a�=��jp�:e��������rKՊ����2!r+����}��,���6�Z4;��M�9Ҿ��{>v�Bi��U�b#�5E�3d~F6М!G#��$�&�����T�e�i��~��%@S�j>'[^�*���ZR,3ǡ����5.\���E� ��?;����̳7������_�����yb�n��?8�����&��	�y�u�ba�=L����o�o��L4*U������I�w5�"�λ��F׬u��0wzAm2�2�PQ!�s�^�a���4�|�y�[�h�R��#Z��L�-/+A�#@.��8�}Hp������?���d�h�Oaen�R�zY�Q�����9�fŸt�8�Q�?�ǆ�xȍ�֡�<�PK+k�4qz��Zr��������<�4ĎP�b��w�D�|u+���n�.5���g�w`�Hm��6Iu`�ghQ\�b�+ѹ��}1�͈y����Ʀ�`"�`4�⤚�#7��գG�ɯ��!�$S��[�.��[�lEmC�Z�$���Ɔ@�<��3�	o|��p��"[+cvyQ�,,i=ǃ��&�u�0�F����gsAc�NKLoJ鐡09�5}�l��cG��ϔ��TL������ܳ�(�u��|����Vs�7$a����5�]7��q��E�"^l��p��kjW:^L�/�0������qj"q���d�:9�!�����H�\RZ4��w��?'�,@�h���>t�z��a̯�9���]�A��>)�5NЇF�t=���i
����
N����J�JYt�h �T0�h0�����y#<�:�4k81uJ��,XY��s$z{4����
żx�>o�@�7����|aY�-�7��@h�^1s8�e1�� t�Á�h8<���5M'}�N���E��!��:ņ$��\N��ZUN~)(���o8$������В��͖��{<�yX���B@[�H�ڄ�y�t�!
D�	Q9}[˘f����Q�L��$K�mMC�R�WǤ�j�Ɖt��\.����;=n�C[��X���b��߇MSmi7�����d��VC�t��;�&u�%H�z ��B	�r�j�hk�""�����4+�5T0�.X���)$ח?`t#
x�?MҀCG|�s
L�E�;����+D�;i5j��~y<oD� ݔ��F'To�T �3�io��3k��	��zY[+:7E!V�����P �}�q�ZU�jpy�щ���-�2t�g����.���m .k�8������4�1�r�ʹI�9'Mf��v�<���DB�2�Bz�����*¡�������z���!�a~qN��-[�c!��ߍ���{�uS�ɕ�L��\z���&-�����ֈY��L�\�i_���9�0��"f���+�Tqx͚�F����}ߓ���'<���#3/��C�I�u!�#�w�i>��\�f���wm׽Q�T��Cg��$�7͜���GF�n�$���쮷�h����ǃA��8=I�C��w��V�-Df��G��+��[ο~���ͷa%[4�:!�@.����^�tû�ӓĽ?�����-�%cIY��xMi�\/�9]K�h��f���Z��3�5��!�R@-5Q�M��RsmB�|�"D�y���L݁ix�B����pO�땐?����p-SD���^t��K�꜄l�f��}rc��N[j�a�Ў11�$�fW��I�d�X>"�(Z
�5�<�U��ҾI$�YC��C=�������	M��H.�e�-����L���!x\]����7]�'o��>��C��}O~�?���'�ڤ�b�&}j�:��U���ُ��l����?<���-�[�w�YHF(�1Zӥ�
��ů����T+�z�w?��� �{l���,r������=��ٚ�I%�Z��p`��*Ӎm��D*5��< R�8��<���X�?-�z�d�NbꥧPJ/�Y���q�#2� ��W�d�8���%R��:���-X^]��'4�
�a�Ý �K��4�����<,y�E��;�X�K��Y� ><�g�C$ދZ˃t���xZL�s��b1�		�D�'O�Rz7ڶ�'j�c!5�09o���'i�	�    IDATO�%�8���k�ƴ�8�3�"��D64��7 �!غoy�u���X+�1�� Q1�3r����l�)���@cm*^7'~��z�כ���6�#����է������0}j�HB~̡P�wL`��]��%��o�Z[-��$�m��Qv-���A�|�ٴp��&3�m�/����ą�����J���\���V`����e���ڻ HD������PЃ���n��� �Yn�-T*ᐦF�^o��_���	��زig�ށ�����>5J~�����[J�<|�(�?��m��(�ش�=}j�}q��@�+M�8q�33j�x���a�]�����0�8t�ZM/R�a����f��in�^T����qyR��/�Aς�h�'�?pzɅ�1�/!�-�FEw��[K�B��ü�<���0{K%EO��܎�ӳ�. /@п��ds%�--�J����(�sP�h��Aڢ�	��b�k�y���I9�⵨j�����CM}�O���H<5��j�Q2.O�kJ�Φ��k5Eժ)bCA�&�rh�7M���"ժ�ժeT9�k7���HX�-S�V��[|Th�ĩ��$���'_��]�^��k�ʎ��{"�s|�*ބ�m��i�+��߳�ea��ǻ<g6�����?(|�hTB����	cں\�~�jd�Y]��>�"��I���+����I^g~V5�B0IY5|�ԩ���ɽ
�.�g
E~VҺ�i��cr"�AW��Bf�dT�����+�?I[H]��"�i<\?4��� d�g�T�;�Ɇdn�q,�]N��'�OW�i�m6fbk�o�/��|�}D�ZH��0���>J��f2m?'u=NG�uE�(�wW֖�b�Q�	5�2��6n��mx�E�c���$K1N�Im5�?R�8,���^��dK��i���g�)mR��d�4�̝���������S�ͦ�T�@���Rw�s����㥃��ǵ��>�A@��m&t���p�^���\���䇱w�vD�^���d.8L�趨!F+D�g�&+N�r͈�K�2L���)���A�!��A�I.Ąe@H���jA������X�6��fC�B%�E�� >�ɏcǎ3���݂�����I��	�u��YN�2z�0p�����<�Epv���h��$�����x�g�q�gQ7@"�g� ،/i�-i�G�Ѭ�0=u�؜���#(�<(׉*�iH��I���tfCĸ�yY�9+ӚU�hB�I��k5��C�!�J�������"�)��(x�VA%�
y�=}�?z�8`����=��o��2L*e0"�@�{T��zn����>��?�ȯB������·��ҁ��D��@fC�i��+jVs8w�v���.F�p�]?��?��NO���[�n�y睏�����G��vp��q�r����%'R"Qn42)����O,����G��\>���U��5�P��b�r/��+W H]���[��ћL�B���UTrk��3��En6���,
��Ȯ��*�K��b����R-"�X�����j�6�oA:WD�B���H�4J�4�8�
U���MU��oaph#�[��4P����7��M� ���;�Q��	�A9x��;�ٲX�����d��C�qP��M���W�@ ���
f^<���<�����!��(Cf:�6, ��Fʐ2ℐ���l�ѷy׼�x�ůE�Q���*ʭ�I�dҫ���cS4����.n�"ޖ��F12ԏ���ka/�aP��<��Ȯ�ėd���5�y�(�'F�;Oe��x��� �����
����M�BؑBϱ�l���`
�HH|�h2��q������
�Y^+�!�"�K8���-H"��)m�lX��4֏���(8|���p��]�������Y/��O~HԶ�۷��s���h��r��r-�2
�
��E���+8~�<(��s���ޝ������D�hz�b���f򘛝�����&�L`����ݡQ7�
���N �@����:"��l�Ǿ�;0<D�9<��G����*���-c�ܶY�o�}�`i9�^:���%M���� @nO>�kK��12��9g��c
��7���*6�Q�3L�� S)� �KDυ�����i�1ב�L�:��W�c<\9��"�$pOS�9���-�zzz�"GytD<ja6*jf8	�:�a?�׫��|�݇b�"��j4���RJ�TC@�G��2�ŃrBȽwnn�j�d�&�|&��¦6Fr [��F����a�T:���'M�H��-��P�T�(��؈�Xt�Z(9�7SkY9�*����YB�*��B��z�D�6���l�l�} ��F�^��X�>���&�����N\(��6z�G��T)�̠7���C%��Ȁ����X���8�y��>YHFb)��E�VK�1	��;�~0��d3�ω�챙d*g2�!KU��j��]��{EL�,�#�Z݊���]�s����tǡΉ� Rg�稵6�,�����}G�E4�41�
��0����!J�4��3��XSf�o�bJ�tS~���2<�ʟ��{��ޥ�r6��`���}:�Y@��V�H*���`�H���Yi��&6#�ߧϕ/�0?;'����(S�qV%���)�8�0��tO=�<�i�39�<3b�}h�`�F�$S	�$��ƶ�Mص{�m�d,2�]ON�I]M��
�=!�I����ԩXZ_(7����9H�П�U��
"� ��FԚ60Đ���AQ��Q{��C��wo�=�?�pT5��!`����0������2�v��x��g104�-['Eu��3Y%	�-�i�M$��-��M�6iҮ�{G��k���LC@tJ4_Q�l��+����oֱcs��w�vZk�:N��JCq��Tj��s��R�_�)��k�ͳ��&����a�8�:�>�� �T;GBc���-��y�%�p]��K�A��F�y�j�<�ٌb��D����n���ϲ�נ��Kg�L�V����Õ��k�|�G�}�[?��cso`�0(�̅�iW�M�ć�w���u
��җ��g�{N�������Ǿ3�Ƶ׼Q�����<�pƖ3�!E���6GP�z��K���T�a5��(j_��� �0��8QTHq�ڤ�� �1�|[(����"�����Ԕ*��t�i��v!?���e,��`��14�VL0�8��p�O�1j̍���^� �;�Õ�)��墧��dڧQl���TC:�D�h�;�bǞ��
EP�3�(&x�Dt�IC�0FZS��X��!P@V�pr�h�)�a��oq��JO�X���x� j�-���P23�������f×�iVT��*'.�"6��n=^`h�V5�.� �fMA�VQC�F�
 9��l��r�%�*�x�it ��:��GctT�H4v���<%�}r�I�;L��W��zӧ�����TO?��<�h��+
��B�!�=��h�E?�99��vn�P*B]>/��6҅��#�,���Mڗ��Vd(!<7N+������@_o�������x�sz$%�VV2J��3�b���c���Pss�k�㒋/@_��F;Y��k���i>�Z
ʛ�Y���G����c϶1��f�U��5��e�o��)�10:�3�ڧ���\#�9r�$��2�79����B�EX�U��=۰{�V��$�=}z/�t��Hb����<1�D2�&�gW�cO���'��GOD�SY�j�XG9�������_����
Ł@>W��\�"6�@�XF��Ǒ�S89�d���vچ{���R0ds�P;#���d��5�)�����*��bU=cr3�S��P�1�����Oaa%?��Q"!:��W'�ǰu�V��p)�
�����9<���ͯ"�@ 3�d���V�@����>l���5=3���9diL������t�����v���}ƭ3S�L�e��B�G�/>�uC�k6�=V�s$*hsc����5dҤİJ��҂��.b�7�-[T�բ+騳KK�9
�Iu���#�c~%��E
���"�<�����d��8�l��̊8豈Ec�M����A?Qܒ�x�N�h�k�Ƥ�����=�{q��I4�2ņ��zE�A����	��"�T���,������x�a�S=ƴ����4(:�"uv�k�M���0�B���-c�-��5�X7-
)���t��y=(WK2"�z�N�P���c�#�t�H�ؓ}�mt�Z�R�x.������RfU&iEa��x):ޅ��CZ+�]�WP�D�~�6b}�<���shx|���D��Wã\���E$�QL� L��ty:��*j8��ľ��B�1E�Ͷ\��8�����"r#r�
1޼y���,�Mk@�i|�d��Kjb�mۆA�VuC{4֟��>�i�3��.KȖ�ZF�͢�B\?��e�p���1&cQq�stn��=?�!IU��'�������Ө�f�ם��F��p�����n��z��N�[n����0:4�5���82<V�֔M�""zDX�p0655��6d�j��{�Msh��5���f�Z섞t.'v7�z�k����s�P6�7/.̩����oG��SϾ��'fQk�4�a���N�Y���q�2�5/Ǻ�)�ʚ��k�����e@�:<�P&N���ɉΰv����K��E40�Y�g���8���h�aW���܊@@�N��Vn���������?�����������Ǿ��#;��;w�?�+���ܳ�7ЛD���,��=��� z��������E��G?����V���A�0~�Cƙ;����^��Wa׮3�wיƻ;JI����1C���O�ŏ:���X�%gX��T
B�M��:h[K5�hŕ��)f�]��&��7�1ݼل�G����U�x<uQi����_Y�@2�x ���9L��
VfO��]E��E�����@�\\�?��/erI2I}�_g�vn�w�K�l��R�I�p��(v���;�D�����$��JNt[
C����0�u�o�y*��D���~y%�'?��4�U�z�QX�`��a����k���nt2�J��~���-�i'�dq��/�M|��w��[~�:�y޹X+�1���L��"U>�6H��27qM�h��&ҏx$�T<��TQ?06ڏDԧ@��y(�gW�92��j	�f��y8m�7�X"�Mze-�����,6�M���/��X/2�&�٬�L�ϥ W�f=�(��܆�۷"��O��k�^)_�ca-���,�L�b~)��7�h��4t�fSB7�/K��5I}k`p8���&01ޏ@��%V�(�Z��V�Ea�o�z�$=�䳢�l�y��32�\f1ST#ݠ���F���k95�k�Ul�2�K.8[ƒz�:L�b	�J�b==��w<:8N��� ۷��̽g���]�y��6�Mo�2+��|u��AH BHhF,��a'6��;�_vv�O�΢I�Fȴ��խ6�ږ�Y齻��n���Rkbc?|P�tuUf�{��y���1a}��U*�O���<���(Vx��e��.�>��o�#�E/I$��8�O��MЇ�zq��$b]Q5x|@QN����*�ϯ�0��!��'�v��az��Go,��G���?Op|.�YzJ�$̻Pk�ƽܼ��2��!�xV&��������m�7��5���	�%}N]��maI�<n��	RM��*޼z��օ��E<�^YJy��������� ����u9Af6���*^|�g��_G ��ˠ#땼B�o�z���jC_'b1���VW�y{�[��4<p��N3�!b)�������f�$&�A���I��^ش����X{;zzz��̴�E��1=���k����mayiM����@ �����p���bC�Tb�h���X�_�����(�X���(bvu��Ϋa�Q�{U$�dWV�T̝=3��[.�RP��rB8L(��F�g��4�W�â�}*o(�h��K��t)��QV&N%�B�hݝQ\�tgO�#�,��/���s�:m6js�˸7�Z�N����(�O�J�3�'>��8ԆF�)��6�I�m�VC�ϭP,�x ]iy�89��NŉC�nAOċ���|�G�䲺���d^OS6e�ff	�6V<�`��f�hpQ��4��)�䆉`n��PK���0iKC�|��nܾ ��=���hs�M�\I@eK�2�	* U��80k���Q܂q�L���cT泔E+%&
�lf�0X���=�]��RX_[F6�ԵB�T"q�?���.93�-T3�r�	�ǩ��̻��悹:ST*H0�Y4@��(��Q�#�ΠQ*i[jmTQ`N@>k|D�fP�Xյwt�^��Ck�����������i��g����2ٶH�~vj���T�(o��ʙ�4�4�����p��n��7	8~��$I�,C+a�<�Z��V�l�f�ͦ�"���R�?ӊ��w���|k[q�͗���w�Q�sJO��������Lp�h�V�b"č�������uS�7���s�5I���q�Nz��"Y<��%btI�UE��{O/��(���GW(7ٔ�����s��ĨZ�չ���S������3J��l����J��+�L�������#�����MO��(�!h!�4����B��B�RF�PB:�eeww���?!���ӟ�c�����yV��'�NN#�L)R\_�E9y����X��V�O?�A�T �\3��#�k6N�i4d1.?H�]�7�49�`a�u���
�Xw�n%�EK�&7�3#�0�^��X�Rhr�%�H�lb{}E�����,�D_��C*l��k�iza=�.��'�x�cxQ�]cm�~Db������,����.�%jr6T���)7�{���5{k���eQ^�|c���v)7�J�������\C�Z>�:J�U�MۭN�2ؙYFb~H�57����2)�\�����_͟�o&�(Cz�4j�ǯ�7q��i�g�j������tRAuMZ�:<�8=!����XG#�]{���
賶Z�(�rҔ�(�_\���v?&Ƨ4��2��Z�/h�������p��֗6tp?��#�SJ"���ں&����Fq��	c��z;#P�O9��&.i;�)l�'������#T����~P?�W�.q�,�jeDڜ?1���^P6[��QΕ������E����0vlH��� y}^\�1��k��N��P/8dB6�w�P�o���d�f�|frO�@$�F�d��Xm�� 򭳽�Qjn����lo �օ�!�zԨ�Sx��Uܸ=�j����Ń>BWW�}�c<H%�(f3e\�~_~���n�??��� �N&)W�g��1�����T�.؜>TI�P���P_�������I	|@.SE�����b6o�4[�v��f���~�ʛ����V��x�����7eG&��Z7zw� &w�h���<��*�-�����+Dwg�j^1�ę�o_����ؽ>8�,L*�
�1:ԯi#ϻt2!���U��9��+��W�Ж���j����uH��O4�\����N��討��ܸy��\� N?j\r2���|7�o�{���Ґ^JitD��XP�16�/�?S��B ғ_�Ϣt�n/�:,.�����X��B(�.��ԉ�ho�p@��(W�DKu8<.dJU�mm��9m��ǎ��1t��(�ٕ���5��%��GQ�rBgP��3�o����S'd�.�/=99N�7�s�S��E&��'[���3�2���RX������"m=��RH�Q��c���(����<�F�`���t�Fg�ω���No߼���u5�@e���6���!p�]�~:,�\Kr��D�E_�������J^�ܔ;�� 6ŷ�R^�V�!�v�!8X[RR1�-�U���
'4aeƟ���?�J�J���B6����hN����kV�4�*�$=1M�L�T�<p��K�a�\
��[M�Y���l�TH;��s�,��    IDATŉb��C">����5�H�����K�l�!�E_;��JF�cH�
U�
W�qq[���(R�|-v>��4��x~F�t9=>��mh8H1��=���dճ)`���2�e�h0B���K[4�acT-��D�#�."�Y|Q-�	y�{��;����1�A���_������/�`�PϢH(�����!�T�\[��a�nZx����5����r���<��#L2�J�^\1�jn<Z��P.s~��:���x=����t�?��.>�g�{_��3�r����v�O���ϧ�G������6@�ϩ[Bz׈6�S�⽨�	G>�$CV��f#�� 
J������	^Ǖ����]��,��dP]��F�A�����J���h ��Q)��ޞ��_{�3�����e�/\�eE��Ȇ�/�����?�BW�����󟳝��jZ�6�	ݳ�(�-"�'ll��4�����D6S�����l��?������1q|\F.�Y}�}��� R5+~��
���Tm1�8]C�P�#։�#5��i�S�\uױזB�D�Q�G���S%���P���!��hj�5��\Es�K�I�XD�i���J�T�z��,�/`mq�tN�;MWҞV�:��s�:��}/*��._�ɳ��׏D���,6��J-�����pƄ��� ���C�!�*&M��o�2��y߰
�ƕ��:zn	l\'3d��>�]�
�r�$����YY�va!���'����j�|C�	��͛��fB�~˸�d"�Yl�
"CC��'>�s�?���!�6֐����uܾ�����vc�hBA/z�06؍�('����m�q�|��^��;w���D080���Ǵ��ح�%_�֭X[�c~~;[;�����sg���&���+kX]����^�CS���A�t�F�)�zN�O�b݊�����po~�IN�c������N�e���;��]eǄE��p���f��p�>ҩ#��G�D�8�$����I�Ӆٹ5��ڛ�h����/���k��.����5M�ؔp�BC;K�t*�����pj|	1Y�l��#ܙ]��^��1�:u
�v?�i������
�:&''0���	d�5ܸ{��.�0QD�N�O�%���x�{C8d��nJ��\��;wp���tG111")��Nb����R��3�g�dC�d8%'�:*8y�S�`t���PW��א��sT��F�g���� F���3��E._��ۗo�q	�
D����h�-cjIŭ�ӄ!=`��|��c�=�a��$@�#���d�@��Prce=�;밺���9�*az��c�2�J�vx�H$,�+�A^�	,�3������m$sd�wj�n��:d[ma���K��?І@�`j��������puh�����&gܬ�p�07�%i��U�Y�g���<��%tF�ȧz���zݚ�Ո��e�u�n�f�g���:��W����	���#� �'��*)���l	 �ˡ��&���0wo�N���sgPB ��p����Y�#�'|H0�V8�� ߏ�N�(�=fQJCe H?�=�K&Ӓ��mJZ�v���L	3��1?����}�1]'�ܑ2{&F�1�ۉ0�]ng��0&K���9�*���`f}��Fn �aj7�_���id�K�KC�7�\�9lfZd�w&a*��І��V'���തDĶ���ZE�eG�׎�YI�P,��Ӣ#U�	�,�%i��l~��aqY����|nz��,�V���Mɡ
s�r���|��&l�67�`܌J1�*�!��rU� L�p!���>*%�ahm�8��7������O~�d�{�f�S(�U�Ѡ���|;��&/�$�7L��
�,��8�in!i�Đ�����F����A�X@��*��5X+ ���jY��);(A�ՉP���n#c1�u#ݡ$�gn¸!(gS���o?�g������5�q����/ൟ��3�������� ����K�Tƭ %]y���C�-BY�P�b�k�e4��������b��6��Mn+ݛ��N�m�^ÓO?�������Ƿ��|�+�h;�/���	��!)�?���|����[��&ZT�}H�FN�;�x��>[a�	����$�)�(���N�,�M���!���Mхa����g�$g��#���(�U�QJ���?RJ���O�ٷ��~�_�����i����Ǿ���}�n�>���_[�>���'����� �.�Z��c؊׍D���_~��'5���x���?{�4z�{�R$k�M��D��\�[x�'K���/�!(��p21��Ҕ[+F�U����g������7�%m �����<��9�2�J�l��N�J�."��"CP�7`�U5�aHH%�j5���*�����wy�=�HJ3��� ¡�X�,��t���(���'�8bL��!7�`���UB+fN�>忓����Zaa�rj�x��f�z�b!�ٮ���kY�f�STԹ�ce��iH�����V�27��a���DJ��.k��j��\x-ِl��Z�bB�!O&���Ga!��}}��G?��O=�d1���u�Kd��-M{-�8?#K�LT�2�GC^�t�K*D?��C�f�I����*~��7��ρ��:�c�;jH$T��Խ���[7fD����(\��a��Eo؍�O�8��]x���w�ڔ�&$�<�#�d����#�_XG"]����TN��Vc�f°L@�}K�]a�����U�ְ4����Q@,Ȣ=�É�R(��s+�~��::p��Yt��! �._���u���1�Ƌ|���E[��σ��Mb�� l�M?���=ܝ[����BC��N���X���9$se��a�#�P����}Xw
�ُ�%�������h}�BA�!*H�������M��GG����#���/�:>�lE����#'H	����@�g����06�	���u}�f��~��,����I�p���泄@ȇ�''1qj��:~��elo��t�t}��+ņ�Ԗٔ4�T\q"RFoOF���"� �B��F�*��vP�r `��;����i"U�W��Yp�X/F{� S�������_������hu=��3��;ʁQ(�|vknJ`�.5ݽQI��a��^�$4�o`~a�lEÖZݦ��𜚦�1[,���V�-�����Ŭ�MadЃ\��<"V��(�8��ʐ�Uʉx�qz��~iyC�c�x�H]60�(ݬ&��,�T��e�,�*�����߾�ޮ^��>��6�κ\��������R�*�V����+���Q�wj���Hk6�,���Y�Ͼ���ϩ�? 9�����p��"
5�HM�Zc�x��菅Q��4]��:�t�XhJ-�\�k���b����aW.����*l6?�.n5��{$i)��f)	F�0�^x�D"���)%i���5�/I ��]1y"|�C��xm�Y�ӆ�Q�k��BJI�J�o��Rg�������HS-�(�0>0n��Ӗ'̜{�	�n� I؞&���=>�H�
�4�%P�N�h�!�|�R��S�!�v���t�u���������oG��ͮgu��':��Us���?��
v䦟�4�PJc+�P^S��X�60�2��HM%=���=7�p�����������bwK��M���r����L�Q� ū+W��Θ�ϖͥӤO�������"J����w��~�_�:q�,.��_�"^��+�X[�$=�cbbB-�A�� D6�l荴��>D

@���2��țB�dʩ���ූQ_�'�C�i�г�8���k�F[{�ȇ�{����������7��Ym��
Ez@x>�"���6�Me���3R�Mӿ`Hqv�\y~J���%l�9P�{���[c�'"tU+������ ����`�tB�}&.���%��x��M�u$Շ�-�.� >k,�����O|���|����~i�ZY��?|�/�ݸ��������'�ddƀ��"�NvH��F��`�����y�[��/~Y���|泸x����)�|tx�PP�!��"ժh8m(Y�(:l�ދ+��．�-��%,�9o�P؇t&!|'/`6��H�`��u����`i"��Q����5x�4f�u_UBF+!JCH�vb
oNL�+����e8,L9��"�ͮT=�*qZ�Ց+du�p��%CNs�0+�����@L]T�o''�l��(k�⪐ &/��F�qS_ɡ2�s�+r��������?��<l&�� drm���*�$y}����f
؞]���"J�kz�_J��ʅ���A[y'�Tg�F�!9�h�Hk����}��XO�}x�=�F�Z�����J���CB���6M�NNA؍T�
/��d�m����h�� �r]�m��O��_��̂��S''��#9d+j(��X^�����51B,���;����G�P���v��P������@�z�([�RA�q�=����T�� ����v�2�7\�X9�3f��x��sj�T���I�H"�{�(��ۈ�Z��ccm�~;ޏ��!D�V(��W�I�ԉ	LN�5 S��*z�9RX�s�;�0o|���N<ya
������,�7/���^�I�mp��	L��9sK��ב]�jas{e�~��mlmH�A��R���>\�x��$������z�6���Li�'��9��cCGgT*�4,.���\�yՆ�����>�:���Y�<1$�>~[�9\������G.�l�>�n�(�J��`���&__���hH��e ��&����dnK>� -ª�Doobr���&��a�����į�m��[3(T��J6�Utw�pz���vd
%�W�74�f�*ϯ���9sFM��AK���>�A�<�=�88-����p
�544��j����t7o�be=�
�r�M0��� )��׭��g���XtB��ݎ��!�>هz��"�B^����El���X������α��Cܝ����&��Gp��C�:��{x$���
R�b]}�8���.*nm�q�˰�\?6���6�~�����*��_���>�6���:1K�-�����ɉNd3>���Y�C^D�^��fNL	v᣽�s��{�,x}�����-H��Ś���E\�����3�ù�����)DCV�y]��d8 ��&�q�{�(��� ˦��*�ݘC:]���#��J�Z��W�)*GM)�M>#u�0ܭ�",t���Xk$�FB$�cS�ϳ��nK��h��_�׆��Y
�@,����P��MA��BF35�w��>�?��Q�l4bi0�jD��K��j���)���v��NO@��i����0o�XD>����$h�k����%��v���TJ�`3O����P�
���9m�4�.Ր�a��$���"�X���!?���}����af�!j�+���Ϗ�˃2�{*P	1� �
2�8�U %U �tk�s�͝��=J�!�C#�
�#D#~����>���T�:�ޯ�|�+��~���E4JUX\v�={�]����h��+M�2�'}��:Ww*�M�MM�9���l~�&м,鰦��A��4����^�I0va��0>���~��(�k���=��~�y�m�T�
�ͤL+'���Uo�b�\{������V)���i�4�V�L���P�H�67�8�<;ʵ����!pZ�Y<�T/7ݽ1���X2؎������i�YɎ~>��,J������>�����_���F�����_|����i.qh����@�/����F?K�͵����ߏK�<�@0����÷��H[>�[���$VW֑<Jall]mQ�䥫x�󋇙Ӎ�ło=7��?���~؜�Zx�[�t�?�U�:0�'�\"�/)I,։��Xx��UhX�Ӧ�I�m�.(=^eN\�nbp�?�|�����!�$pJ�鉌������n��j�}x�P3ȤV���ժ�5I�QѮ4��ć� nL�ltlV�,�M*`��E���7�щ�1�P\�	�G9�a�.<J�x�rE�i���E'r�"��
�X��|KW�a�� ��l�q���0l���jF��������T��CpC ���ߋpg'~�Sx���B�e�F|�\N�o:>T�`c��|��AyL���˻� Z��c��`����v�:b] t���č�E�:ur�>�P�!B"Q����X]�UcKiGԃ��v�u�����pa���ʠ����I<z���c��73�	����pq*ICdX^�cii[�t��T��Ԝ�rZ"��[+F��s�a�KՉJ����p�3�J#�F%�X^�������LNM�P�OK�]��l����eI�
�{�~_���@L$��|��W���Pʧ��Cx��8N��"1���T���Gow/�(6v����/�`?�k��I����~LNG{W�TU[N|���p�<NM����h[4��l2���Awo3�	�w�Gp{\��VGoč�'hp�@��K�zk�o�a+�Ն�Y$^�M"���f��=����m��"����gC��2'���eУ�ѕa�|D	��	��^�v����a��R/1|yI
�eVV��qgukH������ ��;��݁J͊�dF�-q��r�12܏�}}}���b}s_zU���k�#}P@�qܬR6
G
G���p��"���H�Pf��͉
i!�a,TL�^o�lf�#`�����\8;!�%�ɣvwv��0�T�@&����i��S#���!w܂t��0y��C~�}$�n�U�����'N���p�2G��r��R���s�$!�R_�v�3�{	�P��
�١^D�m�S�_��d�<%{{�ً#�+bp�}�AT+LǶ`}s;;I��(o"$��`�fL�O�>��W��R��յ���Ur�k�+���만��],�l	����Ї���'�pvz�7�Vȷ�JTe��ys����	���΁K3��Ŏ)jLc�$�fa����S�5�龦���D�V�!���gM�����PC���`6���m%�Q7O�7�9���Yg��ƃ�s"��E¬5�)��1r4e[/�JW����De��B	�۫�)�f��Xb�R�WK
$�~>�q!t��gF0��ĉ�������6ko�LZ�*C#�ڰooo��`0W8Ԧ)��z[�G�x|�3�Kj�eifJ4ͤ�7ZFt^#�B��8��q���a�3�\�6�?����h�S��9�y��e	���#}͡m�ڜ�{H"b�������O��L������~���+�bee�<}u��< �c�k��:�;$)�5�<"���Z�M����5�5���3�tV�����d୛?ϯI��ֶ`Ʒ�±�Q|�����}����|�Y|�k�����Rɸ��ҡ�%``��Ɛ|�&6)��&[ͨ$D-�s�<��
�c�D8w8*"_�!�LL�c�M%�;���ys��GT�<N��v�6U���M�g6B��m�����������_�5���_�����^��'��z��O�ҩq�}nƴ�4o*�s,Vmv�wv m�������ܝ�������޺yG	�;wcC��sm�$ZP�Rw8P��pX���߿����6��a�=�h4�
��ڬR�(¾��}�@��|&�N�s�O�|�؝�S�{��@g{Tk�%)%�0�ީ���|2�j��DU&�r"C�J�alN���3M����H�k����6ӌi:���a/��p��Z2ׅ�1�36#�y4����-��D��Pi�%}~�gq�ˤ�I%u3��n\G;H%�D�``3��/��X�v�6<H���66	nd�X�����e� k9/�7���A��<��]�@3�J,|�����{Џ��z�8��(;,�9<D*�7Rŗ�K#�knd���l0殪����F����������ԗ^~[�+r��z�!��~JU�88�bs���{��M�@i_gcc}G|Hd�X�����2��I��v�x��i���g�oyu7��Ӵ������"?P�Ģmnn��1CY&��d��=6�${��(��6    IDAT��Z��=c(�����g���ˋH�������iP�i��V6�T���crbB׻M�
�ٌ���p�\+����a�8�mg������ݦ����`c7��^�V6���|���$����Y���]M�'G02ԧ�7��Q/��S��"
Ӟ��XトDB2G�r��kWp���� ���S�>5�4�%P*�5���ch���Hg���},.mbaqE����8?���&7$m�'�꛷p{>��ŧ����R@9��.���4&{A=��<Ә&L~='cSq��o�hѽ��%W�#�3�(�|�ʠ��2����G��簳SD����D���@oPj�-N/�9\�ys󋚸3d���ΝB[$�	^�b�V�s�H&�:�-2�k���"����!iG���faqe+�ԵѢC2�fւi�MC��N~9�Jt�KoC���h�����bVXZ[�R����:� 1@ο05y}���lXt���a/~�p4���^x�V��d
yܺ;���+�t�w���NO��G���2�7v�D1>9����|kIm��ߚ�7�y�sە��k���!�wG�Ig������%�r�:y�F��k�X�XZ������e�M����}z/�-=�z�"4�E��m���Y��"��4�q1L�Xwq��mg�5l4@�jJWgfȩ�S�vA��Tx��2^{�&r�Qjhр��ʴT*\�Y�j
�c��?'��D�kN煫
� 1[�'�8����t��,hCP��F�&C^�f3�b�9eU�z3��5/�̵�:l��ՖD�u���)���_xq��������m$CT��`5S�R�R�b5��-h�	�rf,���_��ӓ�$S��ڔ���P�n2�骻�N�!�D�mh�`�@�_���|�y������@X�5��+`��+���pSρ�H���v����J�<4:��g�<�4r?�G�%�v�e�V ���_C�#Y�Z�)��K�����A�\Ѱ�4��$l4���z��<�^y�4l��2N�;����tOB��&������2���Ď�8�{�@<�G|���!�AWW��	6����z�2�KTl�0E���(�ğ���C�>�ׇg�"���o�ƭY�J�d:a�d�S}�[Z���(�*T5��V��.��2�F뚓쎅���<�(���h�����J�-k�:�+e��Lz��gho���䐚�}meU5�6z�(Rzd3rT�c��J����'~���~�/~�������翈��kW�N�?��������C�N�_��GpfbTd N<-V�M+��T�R7ig�T5�,�3�l�����^�)�z�2|?{�1�����
��|(S;N�É������o,����ى�4�c�A�p�׆�X�V���]��y8�^�Ua��m�ڲ!���.<��Qb_4 ���O���)�|1�:��1W�$�n����L�~?�*$l�`mnJ�7�Z�p�T�=><@ü��C>��pju�*P��p�'���Ѱ�k ��Mg��4�h�̈́�*�_0@�پ�\oQ�X�v�*Cs�������>��-V��9���&
[{(o��!hm8M0�!�!��_���/5�T����~k5&��j���;<�'��^L�;�L��x"�l���XM�śSH9��)�4Jē�Gji��T1趢�͇��>Cm���d����Z��r��'.���g%�� �,ck3�����]~/�F�hj@�= 2��֮��G�I���pf�8�>���7�0�����ɓ'��$�0������,�V��į��^�!�3����:�&��u������h�,�x<h:���FW�=݆��U��������Vd�<q��C��@�Dԕ��-�5�H�9e"4�͵M�8�d`?�C�w�7p���%v񺶠+��vL���������=��:q��iD:���Nf��v�6gWP,�1�é���B�V����e?{�0�׃��zcc�җ�Frr��M����Gpb�\���h6�����W$�ů>v=�n]?̄�����E\���Lن�.R`�	ΠV6Ee'���d<a�4��7������㵬�X�2W���v*+]��B�u'C
�x��)�#�2I�����/!��+L���al��Fb�Eð88�p��],.��~��ڂ��n��԰p������;8�?����H?eE�h�R���t�� .	�7DO� ��+X\���;���;�u��ǉ&�$�H�۔=�Q�\��;�T�IhbM�1�(s�S_o ��+��EogGC�*�3����[;;���bd�_�E^�2��-`u�@��Xg7���b�x?�n��17�$:�"'ϟ���)�H��6�����7�!W�!���Ǡ��NL��O�� ��#��H;���ҥ�8�'�9��4n�^�Q�<�$6A�� �u����qD.�H�#U���'�xH�4�͹<.��x᧯cviVg NoH@nR�b��� ��Ch�h�p��{��Nh��I(�=n���"+�Ԡ�5!��+�t}������R]�&��Ak�X���͢�`wy������*��8�3�N�3��K��-9�f�e>_�y����8=C$~G�c��m�FlprLg�An54��+}�\��h��r�v3�u(���f�
~�Wޅ}���h"u��<�M1���qD�"�������8n���tbo�������o=��e�!�y�P�����j���{�7d�6�k�f�BH��kq{%Tͩ�	+B>�ڸ��R*	{S������@4����Ã���4����ZS��-���?�G����� <VkC�֯~��x�籲���=�yGW�NMk��a*�$�pI�"e0+++j�+����狺~�K��c��l�l�]T��Ә����a�����Y,/.a;����5�/=�?�>���+����n���6ů�'iS&*�ZZ�y<�z"`�E�C�b�(�T��E�UC)kW�M:�-����Y�8��0��k�t���~OX��pr G�%7%{񸨔�YГҬ�4�̱��s(��>���>�������i4��_����+'������x��ⅳS�����}��2j��y��d3P�^��bӃ�:)m��k�y����|�mqo[Qd|h0���F���~/��|�Żx����!���2 ��4�`g{��!�>;�ռ�47���h��cM��!A��:��Y�i�L)N� �j�Qb�ȋ	��f5�Q������`2҉��k���F��@!�	������;��o6���dh:T�z���Hē8`�r�`̵���ʼ!3�4�D���:�:ۢ2R96<��#�u{�S�ce5���m���P!O�ON�x ����H�!>��)CĜ����}���7�C���
~s
g:M�0�����͂��	��G?�c��8(d��L>h��'�����A|`jb�Q��v�TJ$ a����%��#��r�|��uM~�.>wv?|FӢ��Cd�5loe�4�� ��۝�ƺ1:C$ꕌhe�@��s���ՍsS�:6L\�8��"{�(	�׏�X���u]%�Y���J�}xT���)�_#��4h�lX�Ħ��5�a���R�c���!�}��v���D"'��XZ<D�(��tN:���~�	��N�kV(�j44)fS�S�@:�����p'Ƈ��E\cM&♕8f�v��9��z�q[��ab8��'�`o�03����6���8�:�ȣ�102(�7�D�޽uG�}�����$=�� 1dus��y]�3�c�x��:L��raq������ǧ�����������M��g�K�qvb����;
d�e�SY�[����&≼���(7j���W�z��gpX��Ճ�'���2�)fX��͗6 ��>6��FQyv��5��m��=��ް
N�g��bn�@?';[g����=8������%�Wn�`ecK?���@g[ �C���0b���o���[wQ�������8��&`���*#�I`aqV��P$���Sh��JJ��r����D�0	�7���9�x�7�&]��e�&�9��o���դ��&��۽�.���
D��[wxt�x|�K�*N��V�-M,.Vvv��=�F�B���=875�����4��𳷮k�~|z�/�E_wX'Q<Q�ݙ��B3��eI>تe��n�Y�܊˴��c�x�Ho�|˫{x��%�492,�vw�Q+eqzj�ΞBIX֪��ܝӄ��^�I+�i�{	���M����֋�գ�6��ͱU�1S��lUX|p���ho���Rg�tⲞÒA�Q�&K�}�󠶿Y��QMͷIG6������(�T̆`{q?{�@�����hZ��rj@9�/��j@zSf|�!���&@�$$xϞ�t
6�ʺ�ܔ�z@o3L1�3"�3Q��"���+J�H�K�<7��%�k�^��� ����p��Y]W�~5v�C�,X�n��nL�v8<���������G/���4�v�R�ai���2�:4�^�w��𬠜��:����n3%>�a���D������B)��@��A�����#���N�{	2D���j (s)����������tm}_�җ��|��r���zǍ��a>����V-�"||\a�-)/
�s�G��=���3�A�M���V�a-C��0����w�P���kv����X�X��G/�>��9~L����o���޺��"���-��7�AÄ�E�����ͦ�l(Gk���~�\+^�u^l��	��T���R������ZbTK O#�^�يЯņ���=�G2nyy��z"͍~�ԩ�qy�!SM�>���>�̿�%j��/���׿��T.w���㣃���b�S	�&	*��*�-/��?��C#hF�wx�L���X?|!/^��x��˚f<r�a��I�Q03��EZ�-���.���Cf|(;j� @�S%G=�����.� �9�+P+hb��)��S>�5Q� �[md�MK�N��4&�Rfo���ݝ�p�h�����j��2T��W1j��ACfeX,�P�2!�'�I:�6�5�hv�t�J�ԇo8�4%��{E�*W�d��kr�̤�r�gK�)i��cՍ�-�[:�C�'��Ӌ��u�P���c����p�p�- ����چ�A۳+��-²φ �Mؔ
ٸFf����	���_h@�;c!񎇁�hl��"������9����O`����	�'�dx%���V���4�4�.

o\N�؄�Z��3��X_a?������.���b��#~L�Źs'�t�t��s��jC@�e�ZD�-�������j�!�`�8����r|d�����������~��L��/��U���&q��]��m��
��� ��8NW�0mM���kwN��$V9=85>�XԫаX��jI,���-���a���f>F1���twu�\�a/�0J��P8���^�4�)�ΗAgl�7�}�����Y�ŭ{�8̖����������G��<Jbyi��q�ol��3�����a�"fss�����^�'O`r���	��q��,._��U���pb|�U]v�|����O^���*��G��#O*M�����:^z�UMg�O��'?�^����L������\�Y��~/ie���T����0�=J(�������y���Ws�k���)�&�� �z��L##��-Ւ�����
j������"��h�|(S���:�����B�l�W�`ckna�]��j�:8�j׆������z����喧_�*��G��~����~��G��?��.��ͫ����Z����@�\�4���;7ഌ���N75��vEd"�9�cp��]�p��P�+u���Z����{:�(#===���[f���M\�1+
e�>�G:�875���`���ǋ/����m���!��#S(cqyK+����&�Pt1bu��;�q�8GRU�;{"�<�ԣx�l��v�K"8�umV�9��qxs��!��c}x��S����L���.���M$7����֍{H-��b(T��ȋwJޒ:<@����U�����f  ��5�,��57���+*Mj�I1n&�d�M���ޓ�Y9� ��V�+�Ѕ\Vt�؜��O��>l���ML����<0��!6�b�棹9oM[�cA"Z�{�;�̚$�5u��z��4'�V�ߐ���W#�ձAa��`CYʤ���48N�{{:����^���Q��駔���$��b�aDmbc�B�E��[0��5������=�+��		�`�N�*�c�:�RI51
�YP�e���5i�!�U�@X��*Q��9Pc.���B���L��m��I���K��,(T���#mj>3��9n'x�����J!�Z��]���������B�S����/�!�XY��E�?��O��W~���I]�;vL�����5r!� Uj��1[g��M"9��X���to�OT-Q�*��,+�P ��a
�n�B�V�G>���G?b��j5���+��/|�n��~����d�[uM6�!����~�X,FY�rɚ	��n��ٔ6eN��T�[A���fC`��qϞ���a9��<0��t:�`{j6E�g��Db�M�z@D�3�#���[x�K2������o�m�X>�����͂r��`V�Y�y\\�X�9k���Z��^���,�I�������.���?)Z����k2d�C�y��i9����[y���:��9�^څB�#���i��RC�Z�����;{����)�l�,�L�� A�=O�c�Կ��3��&������g�K��ЦL�t⭴҆pw��+̃)���x�.�����2���j��2Q�������s��[7}X��IKvXu��Z�p�K(��+���S$�t��=���:�x����4�6��Ȕp���y�7P˒��!(�f��*L\��U����r^��`y,�h�+f�#O�����)|�����ӓ��88ܓ_�����R�u�6%G�5�|?���)&R7;<�H_D�Q~^�W�ͮ��7/���h|��I<t�$��Je��Nk+"?Qk���ر~�X8ȼ�@2��̝�nn����B,F�0�]�JՆ�˃n8�&=1��h
���+�{wQ�ѻ�FQ�t�� U�W/5E�U۵r)���c�8>܃H�����tևG\����3$1��%i���ѝ�-N>����a�Ϧ������G�rX�a�y�8:�U�-�4劚l���+�'��3�8>ܫ��L��ٹ%M�YE�N`d�8����:�V��$1%!���� z�{u�om����W5M966�_y�1�,`�9=n5���������p+�ukk������
����w=��c(T �Q���x������&7|��$�^1I�E.�!iZis!���(��)!m�Yܐ�e�,fͬ����F���K�pa�S���� bm
�;<�a#^��f�{i���*mC,Ѐ�nA ڃD���._���:�?�����Q~U�P;���y��]� �����W����L3��b{sS�������pe3���}\�YG��LBpF��V{�Y���7�(��
K��Lq���@�ư��6ż�b�mDgg7�,��ҶW�y���`og�Ϟé�,�\B
�����El�;w�ΨO��ҹID�.V��_��{j��Ϝ� ![*��������	�p��$.]8�\��H��z��^��@(�}�x��Q��[y\���{��8��`qF���l�r���0��t}�`�2FR�������YX�U�y}���_� \�����LA�7!V�2�,5���Ņ�鐳2f-�&'�Ҥ71�|�r[��<�[���P�%�� E �����S3�0�hr������Hw;�3x�ߑQ�zzt�Sޣ�>��+���-������$�s�h�\���*�˘���dv�!^?�uE��)@ᚤθ��/���v�	�s��8J�!���    IDAT��yCUv*�����ꔃ�14د GN�w��a��q����>�铓pY��Be*h�V��G�S����ug?��WE���ϠPj�!�k�{��$
�|��߫X������bq
e�r����P�"U���Je�# /����L���S)��2K�p+Iw�h_�e��pJ�
%Vf�^����K�+e����S$s��=�s�H�����5�rK��P3�������`����C��I�VR�Ӊ��#���{nml�!f�̕��0�+��YN�yVpk�Me������n��?�,Ǝ��{A��w�<����)����?�{����n���eά>[y�s���Ys�k"��u��6xn�-pP��g>'�nX�~�C�(��!��\��(]w{%ie�Q�4pV��<�ʥ��3�3!�Y ��oXل;d'Y���MŃُ����~����;����7.~�k���J�~���A�=u�~⒘��2����9'�􂫺F���+�&��_��7��?��᳟�oP�����?UCp顇14ЇZ���~�ˉ�Ӂ��2�}q�]��~Ƌ������o�{�k3o �v��!0]8��N'O��7�F�җ����n�Ԭ�l6M�[���-��ea�cv��hyZ�B!#W_bN�.��������dU�)G�D�7�~�dh���'/f�Ѻ��?;oLfo�А��WC�烝��C��I$ꇤ����7ڍG�z{�G��۰��Bie�p(�l��������7,EԸ���I!Y�|�h"�{����R`��J:�8����|��7QCxt ���`���&���#5C�x3�Vʭ��/�<lLC@+����1�߁��0~j�(���Z����E��x�P�>qbv��G����VV�����g�ctl ����F���x�g�O�pfz������hB��M�.$Q���i�v�YL�^\��[oݖ4)����t�ZF���д9�K� )!p�=�E��a�DP.$�)��}}�7n�aq� �E*H�wQ�0��ax�,h��A^��D,�<'4�E�A�����z����D��A�\A�(���x]2��h�� ���148��� r�f���J��l�*��p��$b��(�����B*��{e`x �h;�.��iܿ7��S$�{��$��:��At+�2�;z�����ۧƀ�{�ܸq�o�F������Ft�3h�����^��x��D��p��d
l(�9�"�8��τ�q���!2�����6��y����bN�m�xj%l33�[Vd�<.���81؏��6-��)�5l䕬�MQ(��g|r�~��`�Lů��6�V�Q���ׁPЇp�'�_{$��n
׮�D&��X��}��P�b�??1���-t��q��q�hf�Z݃�lw㸽�.|)�ԡk:�������w���`������G<w�
������N1���$�x}���҂Օ�ܹ��Յ�g:����7noȀ-iAvѠO=zR>J=���Wp��,� ��O�ы����&���Wqx�����E_oD�$�L_���윶���������N�D	w��p��
�"��n��W�0�.�\zǆ;���itE�!"�-`e'���������=�K�����mtt� U�i�g���0U^����h	���@)�]��g��P=(�U��YE	WU�2�����w��zF��<�!�/s�%�u�>�s����'�03��"1"!�� ��(ﮬ�]yW�l���Z�D�6�H �A&�t�L眫�+�������o��sp�&���������$)�4� 6�d��B6	S%�]=m؜��K���T6�"�G�T59��t<3������jh	x�Ha�q�Iu�i�㸮D�'�J�$�Q������؀�W\���{���]QQ��� nq|Ϯ�.�%$b1��.`yyUt�MM>��岉/���M1��hm��?�a|�GGk�4��P.��މ,���e���୷/alr�H
�
�NZ�k��2Pap�����ň\>)���$�2¬j�hdbG�<�
�^7�^?r#�6\���H-�!��c��f�[,Q6�4�ؖ �����[N�mlP�g�$����#��������㏢�g����˯����FX�����q���U�@YY�۬J̆�����\N�'i��~qi�v(9��ó[�ԙ�d��F���k�^�DJ�5�=�k����Z�����x�/ICƠIRn]���[��qR��E�i�A��9��	��	Ko�Y,Ek(q�[�0�|�wQ5�bE�M��d攃���Y���0P����\Xm���Q�Y-���u�wZ��� ���j�&���Zm�W�(�W�~��7���o���S���"*���=s�O����J�=���g?�	�s�9�x���1�tb��$U�ʎ�q�x�g��+��`~�7��т�.^�i���+�E���*��:T�A�l�ݨ���q��2�7`r�̉�pU��o-`u�=d6oAW����`2%g�EK�'�J]��j�&,��5r�Tl�D��s��&!om�Rc+"'�q��l�{C�Ƣ�]њh��V"'Rq��^�P�U45}���e�e�6��`�O���	/��wUE��=I���LE� �C�:�8t�^��T�,�S���)��p3�cHO� LZ{�*U6[j�Ϡ7^��2���{$��!�[���'���^�F-��O�����%���*�Gn�x���9�����6$��.�]�ū�&�rX�!�Z��w�5n*����&f�W��E6���6�9Y�A��e�9,έcfv��:{:0��ͭX�vAj�70}k�Zw9(�`v�Q��(�ne�Gx1�B5�Ո�������7߼$4.��n@��e6rP�غ�E���?��ݏ`��v8�W���z#csX^��P2�h�˴6����Ƀm۶���H�\PR���P,�B���]"�#ݪT("Z���B0��d��-�N㭷����o�������m�\3��BO�@T�/��n�w@�0C�
1`�8����[�r���V��ъ�'�c�`������)�yҒz��4:r�i�Kh6��bzzV�l*��Nǁ}���֢,4�CE���%�si&g,���j��� ->&�Z�-%(�Y$���ɪ03Bk
8���ϥ	��>X�KR�%��d`�UpYp`h }m2 يg�豴��7��o��k��ۅD8��!�^����e���h�hA��&�Z���-alt\ޛ������D�����i��\��iŎ�n�)�
��B"_��jo\���LQ^/a��H�?ٻT1ǽ�,�yMnW�pq���R��r�\e2�Q,�Žj7�#^�����G��������p�LH�"���[+�dU�W2����{N��]�p�X߈��/HƇ�⒂p��n����K��[3�96%t����y�Q�RK����Ņ5�c9)���8s���nq�47W�7q���"8<m�:=R����WX��éc���䁁��|3KK2�س{�������obv5����U:���|�ZV���
���`1pk*���י�����G��B�d�>H�=�-u^5N&ox<����*dG9j�5yf۔2h���pc�����3��bpx�r��L��T!k��-��iѬFUCeV(13?�BA��h��EA8�q�s_6��j����ӎ{N݁�����h��s�?KL�Z��Y���z�nMH
6��ZZE��47���il�/I�Щ���W�v"��}��6#|�#[[���ūo]��K7�A��ѷ��)���R��m��Ao_;������]��-B+��\3!K#�c���MO���<��px�a���Q�ĐY^�YI����nT}#��	+��S�;J�O�˧���T��日! ]꽋�q��y1���Ht���P8���)��7I��h <lP) ��܌\Q�
R��P��(E���G�Y��<�u��O�C���9��U�188�Ǿ�(�臡�Y����O���t�`Q�R�X�����9)v��K�2u���T7�$F�re����7O��
,N+
d 8=09�(Sd,e�^��l\mn?\� ��*�4L(�0����I��sO�J�g�vlHs���\�8�*哴{�C�������w�)�@�g�Y��|��CO����uƽ�����#�CsqvZ��e^$��L�5���b'�Z�}��O��˯���_|��p:=�t�lpg�>��D�#M�l�	e�Sk%���\�jf����z�uLc��y$7'`�F���v�U�E	5d��q��`j#�yv��h]���lL�����qՌL�E	B�E�{MR��N�Q��h�h��N�&�\���X5K��v��*�E��~u��3�l���FJ�h�Ֆ�'5��T�L��8�}w܋�ˏ�D�bM,�t5�k!��Ca~^�E��SD.��5�<��IR+��W�hI�����6N��4S���MY�B�__�m�`+�BdsC��(�2�=�x�t�PL��$]��5eجftw���aC��+������1<%A&N'7>=��mt��a��I��ı���xr�Rxq*�⛼ϙ�YL�O��pុO`h(�J��X,!���)Z�eQ�Ä��ǌ�i@Z��"H�怛7�ƛ�P����D�^ձ�R�>�Ζ�y��q��^�����r1
yē	ܚ���J�"E�tqK�V����ׅ;�>�kka��,a}m�-ݪQO��=(�fCJ����2:[ZD8f�D�h���022,����.��6�����ʾriy�،F��٠u�E$l�	E��j�rQ�.�7 �ĵ�1����=]m��P���Z�z��A7�r��T2�d&-��r���!��R,z�f�O�U���tt��E�\�H"�w��K�]1����H!��������.��v���O�bbf�RM�E��[d �l"��)W�D��F l4��

�8��<z�8�k�ۚQ-�K尕�ar1�щ� ��:0��mp�)d��R����[X\^A2Mo�\���&x=.���%����� �o�AoW�p�C�-q���H�ak+]9'�\}�$E{�P�Z4��P�\C�b�Ѧ�h��2r��MMD��3MYL�FTJ*=��˚��|��L��S,�����Â��>����=��#�$J4.0�V�R$r�1����u+�zo���v'O�Ǒ�%_cvn�޹�P,'��j�@��w �����$��gj�;��꓀���Yܺ9�R�.�v`��9��ߊ��u3&����a�ce�ݭ��qldԗ��Ρ�Ɇ�G`����N(C�vВ��a9�\�Rei&f7`v����H�Y|��{.K( �.�@ǩ,9��x-e�O$�{��ƹ��XMt5��aPmp���g�& ʗ��}e�,:jHe����hs��ԗ1�
�/�C%�����ڔ�I���h�Ҫ1�â�D�,�*֢��S9
:D{G�YA�qRl��3��M�]�+bQ��O��>(�<_+����3E9��Z~O�É�%���{��	��l�1?7���R�-8,&Is��ÿ��;wI4�<�r��������x���$!wm3�V9�*WE|/�F��w�ß��;��	_�����އ.��\E�E��
��y�u�*�:�"��6P��`u�a�bb�O��RY�w<x�2���<C�7�Q��:��E�yqY��n�����#c��q�/(���$�#l��^�|Y����1#%��������!)��V((:��  f�e4� �l��i���Q��Ҏ�� �j6*2�Q=�+�G
E6�m� >�Gq��\�>��~�:��N�\%-W1l��h(8�cv)m�����QxL$��?l��F����yJ�2jْ�--�9P%���\�;��&�f�V��Sh��X�D9��$2���C|X��%��׃���TII��z�! ���M �č�}�����{�<�3/z�'��nkk۾��U���z�?�H(�|�(�~3E6� �ln�tv��'������g~�v�އ'���bO��ko	z��;���rI:�� �͎������n��Dpv
兛��XG���Bx+co#�:�C0�r.3$��m��#�%2��Z��ps���d#��:���A�����
�1�ol��B��=��F�Oԁ�b��������KWS���|*�N��W�|V=Q��W������&��_ţg�"ŃCw��g>�����h�����bM�͙y$��QK'�3r!P����4ʐ�[U���R��iX��K�n�ZZ#&;Sꑯ�оo'���'�هH&�<=��U�$�U�M-[7���u��K{IN�&�t���σ&���mX[+��w����p
-[Z=ص�GlE봬�G�>�M��P7513�R��M�#���������#�����n�B4����� ����*�M��1���G2Q�+���X<'�Y��)�5��2=���9t}8z`'�:���^�A*����V�["8d@K8��$c^3�̈́`k {���U�9I�[[_���M��D��^�|>yƦ��0;3���6q������`������Qq�ٷcz����"�I7���-lFRB�(�B�f�;���������:�2�2V���0��X���ؿg>�Y>/�G1�z3��Jr/'Wtㄪ�=��-�YR"�-\�r�l
>xv��G*�E�"�R7��q��-����x`6�`�W��s��!��҉z'�}6p��DcI���������}"�n��/
�h�ɘ8�(�p���ۇpp{/�����Y�o�16��x��
�i�����!p��LƢ��A�˫bH��@{��A�\��O�qs|\��L�#���LNnu"� #���+�KF��w��c��7��"�)b#����ElDsbyJ���tsͷ��[ziP���#g��5h��+-��fo@�5E�D�*b�@㝻�I�lwq�X�<���Ui�z%�&�+c|r3s!�*��k�GWlf3~���ɵ�yk.� ��[�[F6�^���-ڇ..�"�N��I_o�4�l��*!m��\�"��'1��b&,��K8��{Hf��CB��|���٘F[���y{�m������ξ��~��sZ�SN�^~�]��/��l��D�F�!�D5P@��sR�:&m��/�7�Et*��9<Pϟ�ݯeH�Q�J(V ���5��ze1��F!l�3/��t�":QC��s%���L�\E&{�ƙ��F�\hA�	�Fb1-����������ɰF�9��=�kK���.kں�BQ-$px�v���>�{O�@2U�&��E��*�t+Kz1�_�wo����g177��	3m��DC(����l=�Ǐb�А�#����B����n�������K#�����J�l�IE�K��]G��;�����KOڪPYLz�*E�&�Qm#�Dg����RO�=�k���jH��x��@<Fm}EQx��Sh����YP���2�:T(�=��L�*⛫h����;2������_��?"���yW�^��6Db�/t[�pTҩ��D�+s.J�V�/�#�^
��7X��b��Y�B�)�|	-�� pc&S����edQt�؉��K(Vu�046>�}d�5�a��TR�nh�a���Nh<Ԫ��D-�A+�c��4�0֊T�=�a����݅�ю2�mRF���v�ZD\��!�*���*� ����r]�LF2��r�-�z�	�%=����ԄR; L�'*�R2z��|�?��_��K���3g�>����w��=_��cf�ۀKo��[#�傳p#�A�X/U���@O{'�9"�~�C<��Y���?�,6'^~�Uy�������@�
ü�Ӟ�\�LHCpc:���U�M6�����$��4zNiJ!��yY�b9J�B�.��j|w)`9�Bܠ����p9�ĆM�?8�W�7�F2��U���q�рjU7�6`�ř��Ȩ�C�f����M����hX6?��j"�@'x\3�M<dH�����    IDAT���(��r`y¢�����߁��rz+��I�M���(f
���_YAfq�XHlG�ey�X\�@A����6�	e�:v��&�*Օ��i��*E�އ{?�1��[��e#��hn#3�.ioݠ_��c�#(�=n�]u��u�`����8��Q�[o_��jL6d~�ӄ�:���P.�a��j
�~�G��뢉Y]Z���^t��y�pi׮�k�D�oS;���A�P��k�Ў!m>c&�w�p�
7t%s1�5�Dw�3:�>l�oE��	N�zI��x6�l�
��)	�L�\�bcmM&2�v�ܵ�U�t���r�������I�A�ˠ(�v���#����ڂ;����6|���(�V��Ϧ��ю` (�D<�G4^kǭxN
x6S�\�8���G!�v�V-���aG:U­[�~����C=���@o>F1�.W���u
�Kkr��s������D�9l6A	ο�6�q�{p��1TJy��� +@Կa5���O��
��������6�f�:��˫�����V\�O,�8!b�/@�xkk��v���Y�Ǵ��2�/#�V}������>x�z���sE̯&pyt�\y*�س�;�Z�9a�ې˗0:2���i�����ıg��m��\���XY[����f�4�������BE��Zhu�&�KD�p�ОAX8�O��܊D�����ά�\W�d�w����ܖn�Ty��5�Y ps�W��:��j���͍���MϨ�T
J�Utt������ x��8bш&c������
nM,"�&g�D��߁�w�۩|�'��q����)�l^����س���o�զ�/���]�i�fn�/��{���[��3h�l�=��c{_�jxL��+���+�Q(�k�&�Z�Hx��*���ýw�`w�h������d������a0�
'���Q\�����8.D����h*�$J��n���$�RD��I9��䂨�v>4�W5�Q�4��k�-�����!�r���$U��f��ʟ�TD�C���.C+cø~���X�����B�SC'�i����~�L$����@~��&hs�|�����h�h�?�C����:j�Nߏ����q��6��]7R���_X�m7�=;��W��ܛobeiQ��Z� ���L"&~�;���g�.	qܿk� ����5�x��7���M"���R7�>��D{f��fh��=�F��݆���/�cy ���W2��ב+D,�s��3]�����$^���q�5,2'���9Ąە��sN�����t6t|dXC���Ei:��,tҋn��ك�����݊���C!�B__��+"��3�lzz�d\v������nw���p���dA1?C#�Q�2?$��*<��gcP3��<�E�`�J ���>�9l�8v�nt�auu7�g�M��%���CO_����sb ȥYQ�DMרb^���ڄ�[7���&���g!�K�}�w���<��^A�4G*��鐡vMg��k#b!L�F�VO�c%69id"!��p����lk�!�U����(&���I��y�vk�����~�#O��O~���O��/��OG����կ}���h��je��-W��>�诛�`��On�/ξ���~]}��?��?n��n���m�A��2�������t�6���g�qm*��)�WCf]�Vj�5��C~q�' ]^&Ŵ�$��vw��6±tJX�����H?,F!�T�7�Yj�kL��G�h�O¡e�*��p��M�͆���}�>$NJs@.&����*���_l7��Y�+!|~�jE�A���B��:u�>�w�8|XO �zv¹6�6YX@au��8��@�S���:��n�	ɗUb���A����EM�TCP���4�P��]�x;IE�7�[ÍV̈n7LQ�̚�֎PK!�-���t����jEk�%��|I���ܸ1�lA'M��u]--x�C�������N%=U�kkE�`���V\Ёc���) ��M%�l z���N ���lm��VK�d��������т�u����Q�契Ի2Fn�ԫz�z��j���ō6?E\F��M�c��u劸C1x�lb&�����WĲ��ptliiq�4�t���&�y4���+66|�,������HDc�mo��m��WO�����O�P)�r:�s{D$�B'����d�,#Z�es)�l���΁��,�0)ۅZŀ�o�7������S��7���"�,2���N��KØ[Z���R�&���b� �k|.�8#qS�|�
&f��w�n�:q:��P@�XA�j���f&�m�������C���L̀�x
k�a��q��'�eL��C"_MH�'��4'c"J&:VB��A=���8�c-^�.�0�����F�W'o��Z���mMp�������Ka������}����8<�`~yM����떄m"�,��069����MI��W*��6��s�rǑ����s+\���L�.��� %%Fkf%┽��`��^1�϶��vt��# ���bcSX]]�����>�@�`7�.ҩff'��f$a�#�.��مMIi^ZY�f
�?��{qp�)\c�f�h�<��p&�Oe���m��8xhP�@Z�2��]��I�/�w�.������C2�ǯ�='�aO�
˴ ����7�C�8��0ۈ.l�TL��1��{�g� ��T��%��ﾍ��5�9s7���h�;>�����]��VX>i��J���"�|n���T?�Q03�$��T:/��D+�F���h���Ҽ	������4R)�!bs�ns��E�4���u=vlF�]���_z�dT��:k.C��kv�U�sV���:��� ! b,�7i�����MJU�-y�]�4#O[���u9<t�	��>�];���G���e��Gi�g�Z3!�͋1�s3��uo���ZB6G)��բCoW;:�mعcN�y�hPx�D97����i���9�L�;��[��S �S*uX-HgR���h6��ѽ���S���ŔL���ᔴZ�x�6l��8�*ƗWP&Bbv�i�����*f����E<� �"Ɋ�B�WT2I���v�㎄v�x��ڱg�v������&�"!����t�ac<K�P�!S�BQ��V%"��N'���uww�����(}�����Jľ�g�\'J�%�ƣр%�8NS��t{]r/,�����h�؍2�&�������>z?���x��7�(�I�\�l��/Ur��FgO;���Ǳk�.<��g��Kg��ʬ+��}�_z�Ӹ�̽�t�m9s�XgP �uD��͙%�t�"F'g��B6_}�b��P�����#���%��R.-hu��,�E�ƅ�x��(��%ԍV$��r9��O~����׮}�����?�Y4l�}�տݹ���/=���+肓3���h%�Å�bE��¨�KM g�%`dl����`8���	�{m%���lV������B�h�dQ�����kӸt+�xՅ:S]Yx����YQM�a���,��of ��e0��<5&�W���-ǹF�1R��i �i�/LU�
SSih���0R��Hl�M��Gm�:�"E>����0X%��f-w�����?V4�	7f1�"�G󿭪	��)[U�����N�l:�r�ފĂ�Όz�&���`�a=�GQB2�bY�����++��B@�nK�!h������dr@�$e���p��!BҌMׂB�6TS0��/K`Uˮ!����ѾoB�-$�����)���̆[��׷a���&+��u��t�t&��ce%$eKK�m^�)��������&����N�͑��l��Y�@�����ꕪ��܁��vi�����7BX]�@._���W���4�~3�M6�#tu��U��L�s���)?��<��±�f
�hm���n�w���$}�zz3Ց(�M�Q�[�h��Lh�nq�ڰ�D��s����y�ZXQ9��k� S�X��13=���1����u`���fifˊk]7D���H8���(,V7bȗj���HhSW�ݢ=��m�欫�`����W�N��@{G'�>�@�V���v��<������bc+_SP���� �ž�;l�K��+8�9w�
�~/N=��}]��E0M4��9��X݌HQ�9p�����@�0���`umC6Tt�`�,��������L��&WW�Y��E�ri�����R�;�FXĲ��zo�7�H"�r-�C��;;��x��Z2�����6¢������1�bfa3��hn	����>�L�B�!98���-�������mª���݇�o� �KвA�+c�����-	ו�H���mi�G�+��2s`A�/���tw5a������Tč����H��d�����n�ua���������{�a{�vx�N��9������-I��7y�G~�mB��|jn	�ˈ$r0�=��ZLla{o3��؁m�ڑ�%����=^D"5�;wW�M!Ь�W��:�2�?u��P-�g\��7&q���SEq5a͌���w����=�r��e�OL�������,x�~�#���f�y>aS����x�Q,ą�`*��ӏ#G����q<Ҹ��.`dt
	R-.��5&����CljZ�H4@��:e��a��A�)bdAKr�r�a�{f}6]�A�ˣ���˿@)�]�,L���m^�����1��f��A��2Ӽ�~͢�הg�8ꅜ��R�&�6[���Z��:��=�Y�w��^���_�|��9�h��!=tc�PI��)�%Z�W%e�`>��tF]��Z�q����ȇZ˴8�y�&~��K����N�#�! �Q�
�v��QCa2��*���g�����H'CJ��z�e�3������x/��:�.�����S�a4���|�*6�4I����P���/
��/��l���Q��J�:J-�Pl�i�]D��\o�$������nh>Q��n� 	⠅��wH��1mH��d���Uz4���ag��	⠆��|N-��b��
�XGF �c���u���:���ƽm���k��Ɩ�lv����5N�s���xᥗ���.<6�l�x6�2I ���A<��7��_9�<�,����^�sF�7�/~�?��[[@?;Je�VK��_�	���X�%�+���R��S���<�}{�bL�0Q��o��:��������� l��J�T����7�Ǐ��4��3G��k�m
�?q�q�y�0��v�D�G�Ɣ8������:=`��g��ML����tvt�;�����p �6W7QȤ���ms(��<T�&�`mr��W.����������%�X�1��?����K�<�p	NZ���EE��/���	�G�&�䬑ʠ�?*X��u���dit9\X���H�@B�)�J$�܇HM����t������:�tg�j�>�Ǆ'Z�x����J4�"�bi�6�a�يp�?K3^#����п՚�aϱ��s��U�!��ą|���f��gf��a�;��-��(�C�����'�,7\q# mIkJ��uecC�
��4~`MMw�FT�u��߅ӿ�t؉X.�͍y_��*�!rT\T����dqjbl�N��H'���\\v�v��+�b���[�[䄑ְ�
s�X)_�h���&'��L9�`� �<9u�Gx+&N�bA��V���f��y-�0��H�łJ���Y��5d`s����*6�t+��2�1#�Dt�e�%�3q*�g9����>���Ď�\FFM=*W�#Y,H����	H&�*V%_���F�'ŝ�붣��S�{\^��4�~�o�^���'��x�*�B>Lx�twv`�A����i	A�j���E�1�/m�6#�(0L6�G6�B�6�u�w6c�@�fz��&��P��6B���ƶ�}r�(J1B���P\Rhg�ezMz���B�B���EO'~Z	��o�ٳ���78��N�ޡq?�e��N��"�FzZ~���Tsj���O���	fE��B3C�迯֧�f��W�II���Ct$+��+��I@_.b���ػMNZ6A��/���/�aqu���#��.7�i�)kޤ7!��ʡDH���KtیD�1�ɢ��Et!�&���+K��1���9�*z�Z��/Ҩ�3h�Zp����lU:��b�rs�!��`�;Q�V%���R�li�LkC��K��rB��8Mع��?<v����8nݜ:'s=}=0����hn�Cx��W��'p׉ؿc� [�Lͬ��ĸdT03���hmn[�T*���ez��Ed�ԗP��ఖp��p��>�3���;�s�Q���B[y��^�2�������#bhҵ��11���pL�CX𲁸��aѼ�	_�X]b��(^�=��u�!|術h
8a��Q�����a0�����&/��ײ��W�r9�
�y�1BC��i�"GPEZ�jnO,�X\�{АB*U-��x��̩@%nUb���'|-'�Be W!�͈N���Y����(��2�c��bM�@.:�4��60�fB~��������C�Q��_�����4A��_�(瑊�@_L����/}�RP?���ɟ<�����1����+% i����f�������u��$$8��Oc��G��{�Q�U� D�Q\|�2^{�_��۶���5�/c)Zq�s��!��kǼ�t^Y�{�.�|�ە�o��C{{+>�ȯ�#g���駟���?`fi3Q|\�.�}���W�l?{�E��/#�B&G-]d6��L��ȵ����Yϐ�]ʉSy�ܻ�oԜ�E����es�$P��/�N�E�ً�ih�4lj�*�%���z�X���h���-��'���H4I)��z�<�'5;���e���Z�Hg2�����燍t�"]֚���"M��Eٓ��?���(�|��x��W����t��B�D2E�,��?���G�����M|�c���k������`bbB8����|�_|��n����I`!ia�LJ�ڐ���Ǫ��j?~�g�r�*�2�N:�'~����	���X6��!�"�sPLOX�n��7.㩟���\IgF����~�
!`0��:��d�����6?�tK�cL�.�Gl(+���;���/\2
�c�����g��ѣ'��/M��8�\V|����bG�7��ׁq%�����"^�0����!���aA	�.3L�(��}	��q��i�A�i:m�
�K+�=W�f�&BU�詅$�N�IC`�0Q�N`T����	dՠ )�&���]%�b�5���U�<1�R�sc��NQ4Ž��t͎M�A� aU8J!@����r#`�b�<E� B�K'e���R��L���c`��:v,� b�:B�,A��'#qD����
��I`��*qA{�>�;(�_xq�P�_��D�WS���!��sEq��>�W��=C�h���*�!���9��r`aɄR��gC�h��v�����M�DƧ&��Rf�N�W�SE��_�@�a	ƣ3�#v�LC�������fz(��t`�S�)���N%�ҙ`�{Ul{5�C�={��kw;��*������2tu�=�A��hj��
XwZ�2Q�%���:�|�\�]~���T"��&�
�f�T����MeU�B��+Z�Z��R)L�,Hx�p��a6Q>�K
�րO,Ը��TTJ%����e��fKrh��+�]r�s��e#0�ӆ��&	��3\�ױ����b�$��Z�sW-N�@h-����2�|���9x�Za4��`RɄX߽s�:}"��Z��!�������N޹�]W��;�t@$����-�#Z� �.���&g������lQ������հ�����&��'yM8��J	�]�8�s ��8�� �T���-�{�&±�tKk���}�K�,���BO��D8��""������Lv;�D(��Q1    IDAT�%�p�S3��p	��1���nx��l��WQ�F�� ��ߋ�N��gRx�Q���(W����-��V:c(K�!��2�*&-������GoO����rzӉ�dP���Ĕ�o�l3��~}Dh��}}8�w/�Z�	����-�gX|q�5xȫ��1���-�hC���t�R�>����}�@�����>llf��ۣ��	�^s��H�e�G{�	��:�ަf�r�3��H�F�(�kiF��/��< Z�`}��.\E$�t�:z�x���1��+M�P2�qLO- N �ʔu�`?v�DS��-:� ��	���a,�D`4 e�Z2��7������~QƢCa�jb/z/��XM��XB&��c�S��V�^�sSx��O�^λ��BGj��(d��I3u���V�2-V�t���5��p��v�w��i )�F�V��b��U��9|��	|㫏�}�"��9T(�����M�ݥ
W>��&�Z�h���H��f��/�^%^c��{��ѷǏ��hP��jvf�?�~�����!����H�e@ų��X��kHg�H�Ҁ���x$YN�������'���<�),NM���ۿ�3�=/Ti��!((�ѱ� ~����о=�55+��#��29�R"�(����F��j��`R�C
�9�$O^�3qo�z�0A�v�Z[��t�����52�����RQ;Y�+��ަ=��QQ�DXÜ�rQ9D�.�<y�F5T�VV�����A+��x����#h
���pK����D6S���Pf��_��8~��x��g��K/au5�l��r��g�q31Գ[8vl~����#�/�q����I�tu��_������n�cy5��naf~Qj("��l.��؇p��	�,��R���E\�x	��v����<��wb�Bɼ�u�O�B"�%��K[g��q�w�zpa"�����+._�Z��rc������ׯ\�ڼҿ�Y(C��|�G/|o=�=h��D���1�PىQ�C(�`*���v;�n��y���F�n}��Ò�ZL�@��]�aW*�'F�~���l�a%��i���8
F?�t�*��&ԓ���22��W�W���h�*=h�0��q�7����S��\��!`�(���E����ȴ�! ��\���)'!� �8�Ҍ��T@�����ZxM�Ŗ�1-��7i	��A�q����s��f�����yHK�49��Y	ɒ���6�>��'�=ІD���L�lQ����b��/,�f)ǒ�{��+�Aq5P��[�#�5��� <Su,��I��*K��?��|�h�Տ�XX��8޶ٓ8ru�a+�`*҂��P(��:���T�!X'߷Z���Ƈ���[��*tU�PU�b#j��E(d61.��5�y5�)��0�M �.�cE���Wk
�b(��TEg�@��#��v9����˂&��ѓ���h=�JbQ�0���f�)czN�.M6�ן���{/mO3E%8���2�g>=�Mf�p�"v����d�)�şѠ�sڳ�q�vv�J��il��D� �t��V��t��0O�h����,(��ً� ~�"����"�
ŲXwwx4��L�K�[3X\Y�����,�F*.Eq�|^�Z��Q ��G1��.��^��dFoK@�C����V�Ji��<,��U�"I�O� ��B,�C,���d��*�ޒ�N� jOQSJ6�s_����F_��u��y�g��]nй�,��M���a��K�u�zc�=Ai��D��r�T�U���iE:15�D&�@��w�BWO��\�F\�x��7��@ǌ��"��lD�@dT,Z��ߍή&�٧B�6:��HR�X:���IB=ӂ�De�p�Չd�r�s��z�]�-��j��N[BR�r���i��&S�B��_��jq�a���mC��	�` n��Y�0x�n��XVqk|k�0
4	7�D#��a���bh�;��Hj9�x����y���0�9���,R���8qtz[�ddݳ���Q�L>qEj��([Y�q�ŀ��0.�{�+[0�Z��3�8z|����0)�fM�
H�2�PJ_y�O{<6INgA\d:y�t�&�|�]ds5��Ai��[N�3(�P��)�69s��{N�=s����N�_�l�	:T�[�/e�}���P����fA�ˌ��-��ܳ@,
��&E3�5��D�Z6��
/Iy�)�Q��ĽN
X���J��#q�1�D�\M=��
�0���h���Oa϶^i2I�I����ٗ��K�`#A�n@2��E�C��':�g�BQ�
"�$k�	Idg���G����q��y.i�I�Nb���~�Y|��G2�Aw� �'���Ь�+O:�t`d�%dIueHu(�3�\g*������~��/byf���{�h����G8����:��v<�_ÑSw#��`an#�cjt��-���1����,z"�L�V�I�
��6���et���D�q�����6�I��|?�_���3K��F���$ϝ��C
5m ���|ѭG���%�jq8U�k����>�|��_��I��l#���XW�|����������e`H}uo.��o����S�>4(���U� e}@��%�-��~����=t/�����_�)��c�у���~>p?���{�^y�"6�	�5,��"�u����ß�N�{
ӳ�x��Wq��w�݊���{�����u��fp��E�{�=�ܼ%N��;y�Їpσ���.,�������λ��ri��~��������q��~��޿��O����q[P7�$�������R�P �"��V�U�4v�\<�;::��x#��V�z�k�|
w�/>�
a�*��B�\G�`@8<��i����5j&��dn+Z��6�0y�U�Cs��"6&7�����}$w���#vu�SԐ ����@6(�վ|J�wr*���	���A	(�R/b�������,�AA8O	��e��>ŉC�����4�{l"$>[�eqſ������Uʤ[ُZ�vI��A��J
��g�a�8�a��K���$r�,6W�XZ�W�T�,:���)-�Л��'͈j䋮&R˾�_�_������7,j�<�ُ�>�q����ŭЦР��6e�*������M�?��� 	l��!W\���|fe��G���3��%	Q�A��Y*ݚȏN\^X��� E��K+.G�E��9�#�|6l�]�]kN��'�MM-�ZhYA�oE�E���:�yoMu �ΠZ��	f��,^�0[l
�����!��i��,`�(����CR���}>�V�Sb^�|Q=?V
���$�۲LԼ�ޭ�{=&:@���Y3"gT�nT(�6�dRE/f��$�%��(��x2#6��r�jE����f�9q/�oBo��M�%�uf�æ��i�4��[=�^Ah�'��q�^���:<Ru�hx�+��'���M�wW6��Ax+�b�"Sy�[��L5��1i��E��3�6I�S�ӈ�
D;�4V����j�Ey~O-EDdJ�3,V:���B�h*y�>��=�r�^�B�����1;��HtK�(F�wv�%؎`['�VW11zS+��雭3;�	5A{u��.��߱�f���cq9�X2�<�w�,��r��^�{�X����B�h�#�c��y��5�]�u���#�$��
��(�8�i��ffV�������&�E:�	�׆�}ؽg �"]G2�6I���R
�n����ˋB�C�4���Ut-ط�W�W&��Lbf�ϕ��.�!$����V+vlkCok��5
���`y $+^J&r���\��lyq��Ǳ������.V��B-A�:��79�`��>b�&x�~��PP%�L�TB��e���WFp����&�����\0[����	�}堅o$�W��R��Ybݍ�u�A��yf����{���1�E��J��f�&�f������$�Ne)٠�ؼZC0؂�;�K����4�Q,0y�H�Ii�$I��J����g#��qF�Ѵ�Bd��Tǝ�w�؁]��Ȧ2�px|r�s��q��A��>�V	�4��<��t0T�8��b1�=���}�Q[[ՐΨ$��xB���z�T��V�=>��A��ģ�	�+�$����B��"<���E��r���7���?�YTsy������߅�탻��X�h��#_�5��013���0'0=:���Q-I�%���Ј��Os�s�Ć���Fs���6�W�̩�Ƽ��%:.j�h��g�_G?��.f4���X'F��:)DH�gP=���f]�F��"��r)�Ώ>�|��ay��f�}Ӫ�t��w/_�w��?���|^?Lz��i�Q<��/��p��qi�~��p�֤��Ya�%-��l�LǏ�Ʒ~�wp��3x�+�����q���9��{_ǃ>(z��^|��s%�$��m��ݔZ�n���ѝw�%�����o�@6���>�1���~V�����?����E�H��*�g��Ϡkh;;�m{��f0�=
˧&�Lf�G>����_R�?��!��#���w�ݫSw9Z�0ڭ(WrR��HW�&���TJ������+Y)�yx0	�����I���=;��O'��G)���@9������.��2<���8wu�L
p1��iF6�(.C��"PKJ(h�E�5D��*-�M%�dQ�H1�&xh���o}%��L^��7_O'�w6��Ft����3`�"��WSŁ���2�{N.X�K�]]���{Ni(��MQR��2I����$\4�^P��r���*b@�L89Q"[.�a�{�=��<��قx�(".�3�$"��������.i��zA	��, ��AqaR�FC�>�
E�^<�T��3<T�pU=X��}8�鏠cϐ�.R�/]Y���>�"��a;�I����z���X�eI'0� ���L&�]"�P!�Ȏ:.u:�"�ͩ���oA�H�G�$>�174���%#`�YTE0����mK_S�6'�,�gM�&베�?�to��q=R�O"i����>�B�8�d}�O8�.r���1�Grڙ�i��W2����U\Y��U�C��(p7�ܨDcC��N#2Y� ��H;p��ؐf8�7��.�Ox$*�C���g���rr�C�Š���A���]�r¦�h���,�;�SRق4�3 �A��#)�D��*��R�u(��4�rU�!&N����t�X��'e��"WB
b�V@PB�`Ӓ�q����Č�i���(kr��FHgd��	zY�aC`"���Ǫ�l"x�X�kQd
�Qۡ3T����^/�����/�&�,$��o�m��]D��B�8�7	����!��!�ɳN��*L�Y���^"��$,�"�.T�5[ܘ�ץ����(6�����4Z8`U�V���c=�[��q�`2Vhr��w"���!u	l
7CId2��l��dfF&��z-���6��4��8�^�3\�6�d.#6�,l���i'�ǜ��y�l�^u�$uc3�յ4�
�[Q,0���X��:��	�-y�o�\�Ju$h���
�`fr�Qح��DC5G</�l6:�x���G_7Z��&o��
9e�ۘR��Fˡ-	mF�&Q%"o�Z��pC+����缑�9��U�C�sC �JKH�kĉ�m���2e�Nb6]m.�N�4��;s�&�Y���Ӿo���l_�]uY�-w���8W��1��IH���$�痄�pr 	� �``���^$[V��UV���w��7���o$��w�9��˗�-��~�y��ۿ� ��",�R�=��CI�RťW^�{�y'�o܀'�|�}��r�"��$�a��j�D�V��Nt�h��x((��穧���U-���a�s#�,�#�AZ��"jk��6Y5�݌r|w�6�|.NH�� Kd��LfE���o��ׯ��2�Wݝ������c'u~�]���ʎc�:+�ƕ�nD�-A$;S�Ht�3�)�����q9�<�w�{ߥ��]/���|��q��Qл����Տoy+�t�m�]X�d��2�siL�C9�-��ȼ�F�a�g��Φ
��Zرc;�m߂ٹI����j�i�g��#��%/�SUS�g���nQ��6@C#���#���csF�O��@�%\���V������lހz��1����I�\�[|&�>����?�^8ѐ�H,aaa����˿�4�]����#���?���������'��Jn
�،�����oy��?��O����ؾ}+>��_�w܂c�f���>���Eݎ��c%_D��S?������������`f�4|��q���� b?^�s������cs�6m��`������#Չp<+�p��f�����{n��g!�;���o=����o/�,X	�Q;�S�D -x��~'{���v�P�\y\K�ZnY~���f�ܱNz�Z� T�A+`#O��_��^>�E3< _l:��ަ
��(��8�za'��/$��a�Ž�D\/��VTz������`#��	`1���CI��(d���7�?w�

c���3Ԁ��Gw+Âa ��"�n]ʍ>S�ؠ�8S�g�r["��,Yl7����^䊶�=w��m���:� /���@V,�T���N�����z�!�R�]9���Դ(C��)�j��QD�F�@#V� ��O|��!j�F]�.���D����������{�6\��7a���X.�^Zԟ�͗����Ռe�h0��M����69r"��CC�����@�����hW)�����<����C��V�?�A�$RGE�37��L��tq�k�6+f[��~��C	�:=�ikZj���h0[=6�>�Q����hM8(��Kژ_�7����)��R�,�.U{*#���Y��Ay�Xx���,�Yf6��9�n8�Z��g]�4�b�i*@�����D/�3o��5��@�`A�2B�PJ�٠����C1`�&����O��bW��5�5P��͜o�Z�Lضy�Լ��!�o�{�:lft(�χE���hX��fiB���z|Q�Z)r��TQ%�ؤۇPb�R4�u�e�h֋Z��Qi��s���D���h��
<�Һ��{s�g�am�+Z w���
�a�7�h
���jF"j��K��B����T�'ت���`2��/%����A�9,M��� �}�HZz�,i5�w�p��&=�r	���P�v0�N���
��9�ZPL#�c��%�k+K��ٙe�Ѱ�.ʤ��DAp.M�Z6|�z	���������T��ߝ��N�aBi�+���YA4��:���PS%݊����J=���o]�l�$Â�؀�/��6�[=Kjn�iY^��2�����WVLNN+�Ո&�X��E�]f�p�$����
�j�8�
)����(��f3n�<��0�פ���(O�%*��dL�}������@PZY�Eu�����U.�k���|��y�V<��K��/|'O����&6�j�܁��aG#��eD��E~N��Ʊ��K��z6�Ә9?j���ֻ�s��t��)"�B��YN�%�O��Ԫ���a."���'Rf�Oa�S���M�OcrrR�i(Q���P.M�fqI�P`�+$���K���^�vѺ�[ai+�f�Pv
�����E\y��(
x��O�[?���et�^���ĺ�硣 ���̯�_�cf|5n�_DH5s�jN�'��̥IA���p�mo����������ߓ-4�wHEL&��H�+/�Q���12I���Ya�MD��"Ƭ�<T���ڪ�/K�H��u���/|��x��G�
�X.��ze'�V�ϩ�����ǃ�x�N��>���Ht�Q�7�~�4�l�7��]|经`zv�2s,��~��"J�)\�c>����w�O�x��G��_Ņ���G~����[���k��?~�GP�P�EQ�5�[�ܴ�?؃    IDAT�¢������\��������.|���C���?�2>���\��*�ƪ�u��l�Y�����!����6��̾w����ȵ�>��'�K��9v����9�y����7�>��|�2���ux@D"���j!�������7�;�߂Z.��-�!�j<���-�/?��s-�b��l8Պ�+]� �A$�M���-�r������&���]����Ã��M1�fڕ �㑘�����^�,A�|i**@����h;<�OW����F$;�$Ŀ���� �J�rQ�RKx�
�$��jf�D�~/�6d̢'�FOf�F�F�H�Q�R�B^/2����7<~,��r����$5��D����,&�Cyn�8�D���lhm^�	n3�i�9������m7-SM2i*�g��=������ʛ����M�V�Ȯ,�����HF��j)�nR�;�u����7h��6�-�]�����?Bj������OG*�zdE�&T�P�l5Wr���,5ޖl/��S��tP30 *@տ�Q%sr[C�9aT&Z�	��{�}�3St�	�ͼ�A2u5_�,y�������ὨU
J�֟%_���p5p�58��
?�&�̈́�������9��<�]uǸ��j��iX�6�����9�Z<0�Ǝ���61���2�7�7��:��A��f�V)�J���/�w��&�t��FL�2�B.����Y4�#	�9ģA5�eMDY@:Tͪ�pR�8��oy�%��2T�J� �kR��U�d���FjŇf i됌N�-*&ݎ?'[d"R�yZ������K�W/jlm�4R=	���+GMן�)z՗K��D�u��C�0?��^�&�����K%c#IosO �~4&����"+�j���I�(�ѩ�� "���U�+@�;�79��Z����0��PY��I�Jut`aiY֤P�H>�-�of.}$_�B7�,�in|� Ʀ���~��`v1)"9ʁ!�Z2��#���F�l�s�����iA[�@V����D'��� b�!���S4�����^i^������:���ޕ`�)�D{��kŌR�6�[��.�HM��p�GGG��m�\?�
�i�h�3��'��ҹ��!��=�Y�\s�Қ���i����p��p�s���gn���Q�I�i�>;tZ��#x�9�"�o�IW���@@ǯM�6�o�}�x�������͛���W~�� �\���"`	٪ɦ��gw��j�Z��Q�@�x�ב��@~y�����2�q�,�lй -S(���`���9� �p����-9������u(��������9Q�]Z'� -q|�9�ynK�@@�c��1���SD���E;�����^y��8�ry<��nL/g��X�����
�;��#g�]�ayf˳�(+��5��@��˯FӤH�5oX���މn��h�|��x��Ȏ��0ؖ���-����<�^�g����Δ����E���]:/tI�=.+z{�e�*������jUsN|����o�	:�q�O#�!�4���8�����?��#��hI���˽�)U�}�7n�����b���x������>f�P.q "�k ��WP�O���Ç?�x˭7��G���
���5���`�ރ�ߟ�J^,�}p�a�h�"3R�BY�B����Ό�vJ��]w�>���~���~���OK��G���y�#�K�#-���*ٽ���}��8xv��/��e�S���ӿ�����ɮ7{:R ���³�*B�e�����D�AH>��X��/���j�,��&��}w܂+�ߊf1?�l�hoǭH(�b���<���W0��b� _��Y��>��~���舲�sW���1��Q�,
l>XM�e��>1���R�ϰ�%��%=)��:mA]ᨉ ��酅��V:4�m0��C>�f{��^bB��5M2����8��T�qs�-�æ�֋��FtC֜��%�j F�PE���m��6�G�g��4�VMf}�|�B����ۏ�҂I�j9J��zk��Y�wؼ��D�ܠsf�;�4�ܴL>+�Ʉ6QCд�ܶ���:����ZI�$�)�Y��60�)�Q(���`T;���Wu��������G�� t�`Z%�<JW���l2���L�	�&�N@t&�AA�{�5x)�m�q��ѬU
���Ó(/� J�6؈����nW�M%���pN��y>)���(�2|�G =�2�s�.u��E���4�d�D)�dR���f������-n��F��t�
��/nQ��ƶJG!
��s��v#�� ��8{ˇr���6���?�6�Q�)*f<����1�RC�Y��J�!�G���6�<��昴lY�#����a$�ğ�&�G�!���Dzl��!�M0C&D�|u�||r�hh2���N�mӔ�TqK$G�6�\��׽f|�9PH���F���*����,�3:SQT��0�%d�M��IX����8�g�ͽqә�1t%L���=#-(�H�"I�%��DQ-��8M�?u!~ګj�!r�B�t�2�RB�d�ƻ��e�T,}~ۼ�u�8�R�c(gy��h�Z�]5�Y�#/j�Ic�P�)Jd��������7�U
�� �~��2�z�j�Ac�h�D�F>��J��VN����o�����/�֘�QU͓^�N�s~�]�.��c���jrP�� L�%g�4R��1�&*�jLc%݅���r6��@�:)Z��Ս�-FUc����G. �Vr�#�.包5���B�F����.����T�F�X��le"-��� ���:,`��a<���b�PH5���6��R^=����Z쭤���s��|����w�i�c��jlY���FXMf
|_��2"ޚB����4lߺ7!�YJÚ�a�u���;��; z�	qcݥ����BKf���f{yæ���ަ)�}gM�3Q#b(�̠�BJ�N�X@��{4*��϶Pp�XX��%��w�}���:�t��� ���cf9�t�.���r��&pjdss�H/d�O�!���<wGW'��D#�\���T��Ƚ�o�Ϋ����jى~�{��'�W>�t��aˏx<*��-(�FL,��[>/�Ѹ�a^S��D4�H<���3J	����M��$(�g"e��E�����{q�[o��5�ܐ�*�zz���gy�*x�'��?���t�Md'�X0*�����m܀����b`�*|���#?x+�<�%.$�{B�(*^F�4�+/;��ɏ���Ɠ�����������Ν���e\y��xn����	5�
*�`�P�YĺD��ɜ֖��&i6��߁�����x�����Ñ�y8M?�%G?�L�4x^r���	s�h�J�Vzf߽������怳��e ��}������<�o�o����P�mį|qՌ����.��/k��pIh�A����K��ý�܄k.ڦ�r*�e��1SbkMT��|��#84�E=����%$-�ZF�I{ <myEQ"��M[��\��BJ�r���E�A�mg�e8�-�F����~�N��4���	`!��M!���X��OD2�|n�R��-�K;��4����i��a�4Dq~��@��t.4�C�� �bLbW6ʌ����͇��ؐ:�@ej�\w$�a
���� ������C�����FDcnRi�l"�m�� /"C��]/y�/-*��V$z��7�cP$5w��Cv����[�2Եi-������m���W�#�%<��8k��4�E�Y@�y�&��D���}�f�����с�M�(o���0`�GII��2����/a��h��6_����E�
�3q���Dl$ƴ�`3xE�����jñ2�
¡����\�����s�g��/�r��w�g܍�l��ś>�L妵^-�Q�[.���d�5j�p�fЖ�����'�^���D��D�q�#��Y�}�EU�������j�Ԕ��7}z����cM]:� �Ґ�]ұ���M���������2r�� �_RY�G� �0)�D��8��b[�]5�VÂq&E�U���� n
e��ƛ��*�"���O�,BFkb���50+	��}j5��wL�B�e���O���7Ä��P�`1�G�
-r���L@	%TK�T���hu)��=#���Mɪ%����"=�iBP1�U���.�բ�il.:G���E�8���"e��9J�o�	�E9��z� :9Z�6�~r�)�� j{�/����Y�Y�09Lb9Yb?U�O�5ekɤ]��J��\�2����N�FAz-_�,��&:�
�����ZS2Z�5}O6�^ݢ�pT3(���:);<t,�0� >�Ǚ L���0�<j�jՊ���`(�H��_��6�%>i?�»�M�~Y��^�nO<~.&F�B�y�hv�1�d��m�U�]a�X�^c`C����ĥ�D��$,&������C5�F8е�uh�Q�~�py��B�I*Wv$�A�c[�J��Zm1�������OV�>w�݂�Q��aZp�RV�%�o��[Dve���,��{�ƚj~NC�j2T�}~�@�"�ڌ���A�BX�u6�w�j��C��2�kg���1��o�SNXv:@]4��ͥ�Y\{�e�붷�K.Eo� j��Ɖ�S�_�tΑ�r6W���2&�g$j����%N(w��Z�hB�H-siW���ǭ�݁ށ~o�M$cx���c?��,Ź�d�O�6�|��٬���4 �����}}}:G�]izD�;u�$fffdMg4"q��m�sV��7N�:�^���|#��ηa��u��Q	����O�Ңv��x��w���x�Ԉ44<�B�޵J�t�e}����OcÆx�����o>�م�B�P����5�[�B��᪝;�@p�U
����;��/�����k��Sϼ���×�o�1���P�逇C��l(M��	oÁ��Cqz
�f�r�����z?��&��{����82�,jhY�[.�嚋1�<=~�|�s�
���{�]�㫿��#?3��~�;���G?�T�m����j�RP�m�e��U��-k��bq�YL�`�A�@P��rp������7`�-h�����6�<��&0�m��?z/�A3؋���Z�ÄU��
q�fD|�yz�k����3�%CC+�~؄�gh����i'G����ni�ς�B�M(�Tf'03���k:I�eG�B(�M4�9&�S7�<�,�W6��@��B{R��M��-���V��S�i"�����)g!�A��1#��Km�4�fkğ���6���&e�NDvA��j����I�=�����N̂�V5�N�̽�/"R꿙&���6畍���t
����q�]��c� ri�K���e5.?&q�g�U9��g�-�(ݢ>�q�����/b���-_(W�Y�Àd�8�	�!���h$���k��w�i���T�<Z!��M��t���-�(Έ�9����CK�#�`�l���Q,�]s��J��͘�`�&���������,��%��-�	l�،r�d1��L	��@��Hػ�M�a�����(ɘ۠8�r�;Ք3p�T����BÁ�0�6���pT�!b�!� ��e&12����y8T�0iZt"e�Pn ���C]
t�j��<:�Pv2
� ��ߢ�ֈ��F�X�D�h��=�������X�5Ի*GhQ���4Dl�j�.���C���#�rCm�����3��
�"-Kt\�-�}Q�x._��<��5Ю]V�u��D���p�OQ�����e��P.ԋ[~�Z�~~n��P���t/>��A�:Ҍ���+Q9 �C��e+��>���{Y�kV�#�e�f��Ơ����U�+�C��;�>j$�`���"�D��Z]BL�ظ���AO�O˧����(�p U"rr�e�f���W�F�M:�ʭ:�#~m��`��f
4 J����?��Q��55k�45�&�rAx<uR|Ҁ�}5����Hq9�:��zC���:�BЌ����l��=.����k��eRp�DʀY��9�^��H����	��#*��[�Zfx��0����ni8faq�`t&�\�_=��z蘁 ¡���hP�d�G���sOʊ:	��s����-2jR�ye��d��J$4��+G��{6P��h!�%-c[�T
�䳨2JՎ�\+ �]@��Aw7֬Y����lX�w>��$�P��,l� t.��6�tv	�6����YR���~�w����Z� ��|FAD��6�A��p��-x��������r0x><|Ͻ�'��`��D�Ğ��|���RA)�o/ay���u���VQ�=6-�cA�^�+w�$Y���شa/�z�<�(B4X��j��V��"U�b�f�D�Y:4���r@�(Ut��H�3�������I�\V���Eijj���{ϻp��;���%D��ċ���{.�l�>s?����].�����������̧�oz�8v���_�SϿ�R��b�_+ m[>����8������ÖM�x������F�'���я�]q9�۽����Tn"[k�iZ�X	����0/�,P�
W)�W-��4�`���{'���7��#O����(��X)�3��홅�q�F';�A�P�|n��,-���{o���|������o��7���|���D�M����oӈ��_f��IA�om����1Y�ZD�U��7�o��m݈f!��y6�I�h��򂡧ˎ���~<�w�� |�N����-
%-����;̦҆����[>��_�L5Ww P�:�F�NN�o�P&��.2���q���.'�&�X�E���\mDCQ}/B�,��S�E]l���T��X.����$�L�ж��>,:Ylk乚	�nֶ'��6H��IS���Dű��%7k�>�!#������;5����&y�Z!�����5��G^�g��@��B)�m1�,Z�h��4�����;oEt��ˋpʴ�d!w��\�d��������S�\q*x�Q�{�}(U�5j�g\Y)aa1�f�R�'n�I7����>���[JD�G8L{�rYK+yC�� j���203}����.�� �E����%,,eP�q�ِ��[.#?=�_�9����"���������V�Nߠ���3�eɿg2uM�Rt�6�8�X��+�'���'%(}aa	�|	�B�b�\A�|n�
p�%B����ۍ�N��ְ�N�{�g4���>і���p�@�vlb�ό���y,���v�.�%�?@
�^��7�@�A�
*	���Cޠ-�B&+���r�=�j8eb��j���ry];�ъvh�+!��[/������p�Mݦ5��m�[�е�L�m_�\TN�Xmږ��,�D!jB,dO� kۚ�H4 ��=�_�(fs�ؖ�RY�)�P�旃�Ϙ�CG"rQIǐ��I�B.��,��C��?3+������3��q�i���|YK�Vԥb
�(5ԇ��!<҈��� ��aN&�]��H� IHȡ�KA�P!�Z���	�}��WZ��!�M�(c?*�*JԼ��6��2��K 9��U3�i�����49��iRg6�<_�t�i&�^R68fK+�����:æ�K%:�q����uBD̟��1�"6u�K�N�6F�//��P/D4Q�*�C���j�Ԁ��'� ����@�f��?g_�@�o�Wa��u��1p-BWď�SG����0:�s�g�J-�(�e3�e�h�^�C!��v4�`<�2�txF+�� JZ"��RK>٧��7GzGN�C�A�2����R~����Im�
�2��-�4h"�Ƕ�Zϔ��@T� f�5蜡��A�I�	�!���}874U����s�e�]K����	������{��N$�](ׁ�{^�W��6�B���8����Ơ���9\���&U]a��뇰z�Q�:�f�n�:�ؾ��R��    IDAT�O=��DXZ�r1�r!+����Un���'E�=P��ש�҂fa���8 R�H����0����,M7m^�o��0��X�zz{�$��".����!�aai�_~	�Sҗ,�s�aE#t��C����	�s��ճ=���k=��GN`a>�/n����x�ݷ���CCC���{?����?ę�q\��J|��~W\u�{�����#fV�(4�f ������p�%��o{eO��|��hd�x�]���>� =�_�֏�\
�P%jO��J�"Hi�;��,��"M7W��w�w�-��3����|ᖯ|��ϕ}�5v� �,���A��6B@�(�y>��<��Ig�� %����c���͸��mRg�5َ�AَV=X,��#{�̾Q����l�`�!Z*u���P�0�V�g�6|^�f��9Y���)BԻ���,ѫ^"M�|,�,�����Nӎ�'i
A���Uٜ1����P���k)tS���QY��ӛP6!0�l��\��\�1��AY��)6� �� ��F�/&�K�R�)�B;̀�CE�qE��^�M
6��J�%ߘ7v)(����/a��)̝>���	%c�����n��g�鹁@��V��@ ~�ִ�QI�;!��7�}�k�1�8�M�,E]t��1��3ĨPT��M6Y�*��tD��G2F(l	=bS���	`y��ӣ3�d!"�0|�:��X��)n�yH0y����<���dJ��[<I=
�5�,�R?�{��ۋ�nF��G0�U����
&g�w�+���M�6�!8k���I6�-#(�@��Md9/>.��"�t�I��G&159�期?[�"c�@��ukz�Q{��_(4P,;J��gZXZRW����lQ�;:��NX>5[6?|�l&y{��'�(���c۶��������!��`�c8~jT�.��b�Sw!����6��� ��*��
Oc��IubU_��z��5,�������	�"�a5��I0K�'�x|H&btm��I�Drx͹��a��,�.�X������*"��i�I�!o[� sJ��i��n; �nZ77�R���3FgGTHd�X�[�R�A$�a��nxP����M�\A*GwW�6�E��J��ȸ��4�
!�~���S
 [���Ɲt/�N�Ye�':
i�`-!��6�"ǥ
��&�\�,�0uGB@C�2�X��TK�����{ܐF���a���A�ؗq�a!DM��Bht&��7"q~)deJ8jw�p*���e&h��kk��%�Q�bFN��@�e�%��b���s��5)���f�^�	��>+��z��IdJ�M��l�	��%�d)f��z�����]T	]�3��hK���P�H���t�PO)
�&�K"�58Б�Ntܧ�h���p+�!�æ�H��<'�� B\'<c�a��Y6���L,�MY�&m/RA/�'G������tg�I��cQU_{- h�����`�d�PK�:w�����/j U$M�ҋ��r u�P+"!z���8��ˮ�.Y7�Y7�5�|��;�^��	���@`�_s����n`i�>�kt���h�����>g���j��`Uj�P,�1?;�����?��~t��}�K��S�Y�9pT6�t��3�3��
RC�i�U���t��'���up�uo����p���z��z�{6m\�M���=8��n$�ADI	-d�-zH.rD"H�#Zh����NkU>��A�<)��Ւ�.����m�ؘ׆�3�����r6ڰaz�Rj����γx��4�#�H"��ʋ��9�;���rZ��y�%&=�U^��E(�}�z�s߻qх�05��3�?��=���>��Uwg
w��v���wc��a+�y|��G�/����p��;����5\�����գ���g;3�\�!�{�g���LGK� �ݛҲ8Ш)c�����;n�'~���<��c/����m�e������1E�V��斅�F:;d��EU��w|���w�v�o�Li~�����=�����UV�yN�l�m&��� ����R|^�#N�ⒺQ�;9l��{�o��RX��J�<�=��kY���[ �����)-+j��-����=R����p��:�hjN�\�a��	���;%�W���@�X�2� ʹ�M�����b�B+��X���S.鰩)��� ړF��$������G8�@,�B<��(�m6e+�
�̀6ܸ�^�l��cN�NM6���:[r>��q�|�k+A�4�<̔�C��,���������'1u�Z�
�bJ��u�]JԠ�_�K0A8<b�ρ��4IŦ��� tN��Pۏ�;/��o��ս83?#M����4� �~ �����h�MD��6�BWR�������Ё#GO)|J��V�0�����;�f�$�)D�aD�@���
r9���`l|
s��j�9TPP�ᗗ#� ��D�N���B_��l�@��B��9�M���^D�v�?} �m,� ���RU���SDg<��kp�%c�'��癜���ѓ���UBAu*�Ė��~x-�QK�\:����Ĉn��"W(��ֱ��"��7թ�c�@�1Z^fHj6K&����C�O��СCr�ڴy#���da�XX^)��Gq��8���B�J� R�'�cx��V��[Y*adt����^��|��Fw�Wԫ��<}�YLL-�����[ab�;Q��TJ(9i�/:�<D�6*��{�vu7A
�9�zQ(8�dȮ0!3�Ņe��@$�D4�� �Ŏ�<�N��=�Fn4
adc��C�"9Ф �wJ��{{;0��_M=�GGgpjt��_��6�@6��H�����:�qY�+lByƧf12>��SG��O��
�m&)d�N
�������m(%�1���B)c�mn�xІ�� I���@(�����@ 5\�n��6_�%��V�D+R�'��v2�R>��:hy�.8⢋&����:��4*ED��6�Xɮ耎$�BMrقI����SB�b��H��!Fa;*����WS`\*�I�F��8M4�M�i5��xL��Z�P���^^���3Pdˁ?�蔃��l�is�4bkj�b���i�[O�ZꏂZ"��6���5�(:�=б�Q��c�-�(����U�Dr 3'`{�M��Y7?�<iF�En�A��r1ۏ*��'��'���8G�]Kх,jZh�`6�DUxﭐ�$�l��5S�`�DEj�d�{	�kDݘ��d�N1�q�K���V����A��2�b]})Q����0k�hl�"h��B�
��@k��3HM�ԡ=�7 B�R���C�;����9�!I�]��6S�qD���-��b)�\nK�sz���^|�T/İ��q��}
/�rDBu!B���!{$�P@]��I:�;|�֭�e�\��`߫�g�^7�%w�u�W���W1v�B4�`ѬWt�)���鍾�l1y�s��AW�k�k������\��@����h�P��B6�F�RVƃ�j5�K�Sd�[�?��ՇF��L�����R>+�l�y:�L虛��G�qp���y���`f~���2�~���7�[nƎ;t���x��]x�'�������V|�����{�u����W��M�����/�na�~Y/8�_|ť���+�th��:t�j���V��/�_K�]/���}��p��8���S�mY۲3\I/ ֑���.D�V�����,V��Үw�r���^��������EŭV�����̝���K�A�g0�هۈP)���ف���QO@��(��ڜk��f1�u}=x��7�査aN�6��s�����Ș�ރ}��� ���^��"�c��n849{�Zh��p!8ׅu���6�j�9y�p�d���(��^�(�w�p2�*(e�1sf�'��Y-�UuТ�Z�d�.D-�7]�n6�Ąe��ۂ�v�`�d
����n�t��G>,,�ZA��Wu�ׅ�6�2�����jk(�fڷZ��`Z�q�ǈo����^�?�ܖx���p�yQ��>�����a���h���Pk�S��i��t��k���p���4ˇ;/��~;��@��.1�;�Oh²<(���!ҙ(�ꊪ�*���z�"SG$dÒ�;s3���"zc�3��D�66�Ī�x=55��H�@P\T�QT1�аTffVpz|JA(l�I��cB�^r��L��דĪ�P�G$�T��
896�#jtHu!�l���T��rų���6���l��U��X?D˽$��{�Z�PǑc'p��i8��z�fh5�ߺ�D�BY�U��ss3�}ʲ2�G&�G&�hzfN"�������硧�S(ii���q���SiG��c(��oڸ������:<���z\�m(�B�it�-��D��!�t'u�
�&N�k'O!�Oc��\z�6�R��5�+��~�;1�F�BG�_��|��U*g1;7�5�{������N��%	��In�}B�r�U�e8e�b{����+�*ہ)T��a.���vp���c @퇱5$��6�`¶]�8�z;�ۓ@���E�U��-���I���"�! G��΄�p�'�]�^8��T���]crcSS�n�{��O��������k��N��+���*kl�����$��$�c&���Pn�1�\��^G`j��djwH25ե�ᗕ��{���Tu8\)ע���Hؒ��;e�IW`o[�V%���_R�u�/`˸�Q��+ ==	D��T��Gb(�+�����bZ]��V�F_o7l���,�FƐ^)"M"��@�b�QA"ɍ���p)6��"���uY�n=]j��l�3S�a�5�#��0:1�z3�p�[(�'Qn��NsE�� �<��#';l2gHK�A�C��N���ӣpJ"�&}Kj9�5���=H��:#�����c4Y��p@p���ցH��D�2��ao	O�������(j4�#�B8�U)�K�-n�#A�����b�b�J�n����Po����	����w�B	
b����᥎��0uAoC��R!�5ëq��m�D�>�1�5�f�>�p��À�ؚ>����.�� }�@C��\5x}?v�"t6��]H2_��y�PH�<�r�dV��i�w�u��}J?�[Q8�����
�_:([��}>[��D���	ѫ`8�?�%g�Htubpx���.-`rbJv�<W6�J�׃S�cf��ৣ���'D!X�NW�lQ��効�V��'b����@�z�N���I�V��-����A���2wD��y��g��s�E����kW��\j��!��	�oP�/{Z/���ȯd���q�v�u�]���/�r1/����g����L�si<�����/�����\vmX����_��o��r/��2~��sx~��/�-#)mA�l�]�x���LL���//>�,<�v� ��O`hU7f�s���?���4F�g�J����5�ᵃ�꺫���+���	|���199^�6�/�s�M�������@����w=�Ȯ�x"���^��1@�=��L:7�� ��4�Q��p.ں�i���S�֡A��-7�k/FPj��W5��Uiz���p�t�y�0^�(HT�@D�J#%4(�~cIȁ 0[Q�x(kc���;�b*��%$N�-�/�Y��΄����)L�����$��4j�,*�����`��c�Í !d�J��0M99�2�� `����΀|�G�\�[�n���mH#o0�"�a��҉����x��)m�kHkІ�+���`hqI?gn�0�5���z��!T�E̎�c��a��T̆Bn꺿D=���ꢢi(��|bQ��O�O��qI���p�%��;���ITJ���SuhY+R��z����-Zs���BG<���B*Aog�3+����o�`���~��8�ɉ9]S�P��:����S6�������$��4�׬���0<���%�.����Q��|�x8�d<��x�h]���I��a��40=���㣘�YA�gÎ��?�����m0Z�s����<Ş�p ����w�+���:\����UN�����Ǳ���`2��/<[7�G���%�܌151��L�"R��YA&���1m��o=lێD"�r�dj��/,��l"M��^^&�jN�(�Х�\�Ճ}������#�xn�>,,�M��gŤ��&����\p�FD�(�y���9=�m��P/6nP�1_#:�U~���Fg�-�2����7P.�Q(,��wಋv�+�Sl����=���KC&�a9� ����ML��a�L�@��>����(��w f����DZ{61>��vaxu?��b���HA1��&3x��=XX� ޑ@ �A"D_g�09MTOg�P(~�rE�o��pt|�����B�����Hz� ���U�X?<��Ta�8������Q���2����"�P��c���� ��]����2��P"����7'H?K%��yzz;��L"�#����+�B����E��,abr�tQt�x8���.l���ߨ��Pw��0���4������2
�_t>�nR~Mz!����O�o���wu=%��cy14؍�֯AG,���<p 5���l���5z�X�I� J�{M;�Bcc8=6�ӣ9�|1Q�X���U���q�A�=�V���/�@o
����p�u�:{����0��v����<B���nXv\��%��x���1+���)sO��y��U�Ap@r�1��6J`����zV�q�l�QO��WX���UHόc�]H�0lͯ��L����׃˯���l�����Ǧ�P����]t�����scC�_z��J����ڪ*t�/�4<��6�l8B�׮[��
��=%�V*6�h�msho��0��ҩ-*n�}�kƳS��m�k�����=<��wQ���e�B�s�.�:��˩��1O�,�;Չ�n����^tu�ѓ�ç>�7xa�^-���	�H?�.�s7��z�fCC�Qt
�Ӗ<�B F3�G3hK�H�����mވ�D�ęcG�t򰘐m��;m����95a���:U!�����f�H[i���:�y�>�}�|A���cD��h���N��(��@�pW:5�4D���\޻JC,〟YU&��	�LV��A�;�y�V�҇އ�n�ytt�Uo�ʒb��+���_�?~c�SȤK��g2K�ǃx�}w�������w�����/��3�:+��zzq��nĥW^�T��k3���?}�>�Y����>��o�>���3x�ɧ���]�	�d�50Џ믻��p#�~��Q|������Ѫ��;o��/�gh x�_~�·�糯�����M9EFm�m�_�ӫ׈C��z��B5\�e#�鍸�����A�:�c��4[�8~]�����lU
u�I�/��������
Yqm���&X�I�R�'��q�}�\E�Q��a�p �VS#8|`�O*9�^6�J�:�p�0��H��\x9��U ���Ь���->y���gg�j�jh�יB��k�]�U�!�٣�+��]_��->:_R�d�H�R��������k@�a��b�*d#�4�OI޼>D�1��z�"�Lc��a���.��@��s��sC�O*���4�OQ�8LP�@�:ۋW].ʐ�׉SS�
a��!E�J%��P\G;Yc�bM�ذѨ_A_*�ޮ��R��Zu.�0=�����6�Bvc�A�ZՉd����Ï`��#��66mތM[�#��%��l�QA���G.Wҵ�DЛJ�� DwW�	~=n��p�^�/�5�,���3��Β�O[$�zV�i�s��J�$�ѝ�chu�!4ky��)p���S6��O�b|v�D;�މu����An%�l:��S�鑓�
�aӦMHu�D{��`߁�
�"�h��M*�m�|ay	�3jp�r��h�­�	�k��7\�����$�QL�-��16��N��TPY��6m���;���g�]� ���ɓ��oٲ��q4y��F�T����bj6���,�u�	=j�|���o5p�[n�@�h |����0�~��    IDAT�/�1�m��]�����v�=�eo+�To��R��wW!u# 3��|��eF^)�)��Յ4��?���R���9�j��BAds�ɑE<����+Hv&�}�H�����n�@%�Qt��zF��QA �z�62�]/��|Fn(��}1uV��j����X���(�����,�y�%LN.k��1�ϢE.�	�;���&��p0�)SS�Ng���\��t�)SoÇ��w�ƪ�nl�5!�� ����8�B��L���:�9����h�A����1����,�<J�Ä� k?���>�b%�K.��\2,*���˻�b����5C�$�d:@G!�[GW2���å�� ��ػ��;.؆���x�l~�p�ŒZR�e�"�f�b'N�`9M��q�[�G&��J��ZY!_�Y6���ѰGׁ��b�A��A(D.�ǩS�p��&�g��'�z�z��NIbM��h�{�q*c항��@R0�B�E��v���TIϨ(�5��_�ci�8�B^���~���~����
Q��t�� /@п֑�i�Cظyn��-���K����� �R� ���Yg,RǪD�~�{j�E2"B��=h�:Z.]5���L"m��CCk�&�mf1@y�Q7I���g�G[n�l�\�!�8c��z��1�omj�����'W0����sLց;��:SW"��A�Xw������;��@�j���"���g���/��498q�~Fu���f�:"6�=\љ0F� ��>,����Ɵ�}R�A$�r�#���C�(<�"hzV�"3�M���0@jڋ�R�$��� c���F��K���L</���2�y�X ��a����@��5�F.�R�D��>�!6`+{���*h��'��1�3�/aq~I�zL�E�Y�x������_5�IF4
 f��x���؏���c��<B�s��Q��q�.�{�{'�t��!ly0�/�����tx��W��{��M��T��v_�ڷ���ݨ�*B����k�g���hg<1���N�F��T�!��`�.8�)L.7����;�>�c'OU����w�~ӯ|���u�ݸ�����A����������w��#҉�T��h\o�D��M#��6=��%����Ӕ]g�� a[ظ����\}�H�Z�&K��]oT�-UQl�X)���{�V���� wڿ	frc�h�&*:��6ȌZո���q�K�V��b�:m`U���>d�ǰ���171���ÎT��1M��iB�\�(�e(h�)���ᚠ2) AmVX��%�kx�&5C�&ov�Z�S�X�z=�_t9����m��һ�EaG�ߺ�rr����,�l\�rR��룭��pW���vt��k(��J��I���e!��ǃ���s�J�Bn��9����8(�Ȁ$
SQzh�X�r͕x��o��ߍ��Y�
e��ܐ�Ӭ{��� Ű*Y�z ��򠳓� 6�bU�V� }����E�-fP�02��W��w��k�4�uG��Sa{���|j�E�XH��u�ѩ������9|�)(Ys���}_bazR	���tߵM�z�/50zf'Ʀe/���k�>�H�a3��X��QUB�[WW����J�Ь�Q)��҉�?�ۇ�?��<N����F�`͵�V˹�U���/`��&�Ǆ��R�����~�*��J����XZZ���شa���|�X�_ye/N�%��DJ�(�Y$�~w����L!�+v�6�8ufϿx��I{���Q�p��q�CB�?3��S�XZ(b�*�O�1��v��54@���brz��ڏ\�Q��F��F}\݅m[7 ��XY^Μ9���qN<� �ǚ�==�(���$:��L��q��}�Ɗ����Ӡ�Z/�Rq��-B>�a?ГJb��]Q�|V�6�.L�022��Oc9C?z?J6x��-l\Ӈ�ke-k�~_Yѻ�C��W�Z��bS��B��_bp�e���Aф�����"
�!��P(�R��K���{��DO��ִ��6(JeC�dN:��-r�2nE�K�ɢm���>7�46`sDKf�oD�ZUXؼi֭�Ҷ:ҙ򅌆�h"
��]���/�3g���}�狸�������|("��r�̲���C�e�������'���p�5�chh����E_=xL�=�o����O������	\�c#���=ur���f���#Ea%y�&?���Ť"!R�h����'��ɩiL�M�\ɣ�ʡ�/�[�|R�8�BU��"�)�E�@с�1C�9u���r�OΠ�z�mv�4*^s25&�g��7��1��M*��jp�>]+	����֜��J6#W�hЇjf+�'0�
��~�#ز6�}������+�~�idV��.s��$֭��o��\v)�y~>��@�PC(�)�>w�sa�g�!�H��@���h�ׄm�o��1�����8�z@Kj
�����������`me?��ݭ�@�X9�H�m�����#jn�������"x�Mb��4��ɍJ�*CO�ז�MC�~���]w��|׽H��K�����/�'�y���YVv(�)H>��Ss̥#u?v4�@$��&����M~S?���U~`�1�z�P #�bi|4\��9ixd�*P.�,�ݶ(f�A�����4Al����U�6�˩.�b/b�]���+�́��R��(}�

��EͤO��y�P,"_*��g �V@���G��[P�����Eh�+�`���p��oEgwƧ��k��x��gq��	Tk������ �_@8���;/�G~�Wq�e	k��5_��$A�i4J<qf�����O<��^��w��jo���{p���`x(��������#8��ޱM[X�a���}�����d�Y����=w���~�?IŤ��W�|�W���������ݶ�'X�:r2���zx(L1�pqֹA��^A"hc��a\�e8�0�a��s�`bi9�K�cH����gO�ɗNb�D�����!=A���`�⹁������a�ZC�n��N���v �C+�H�豁X�����8��Ә>y(�h���2t?�V>�
�!�� �cnI
7ZH�:M��n#�X4�C(�9&T�ƥ��Q�;J�<A�H�v\��;���F��G��@�1օ^+$G�S������d�Ñ����
WC kFZ\�.E~�_�KX�����(�͡��{�`Y��Jou�9�нsN'GD� D� )�$��#���l�l_L�/\e�G㱲,��� �� @"���sv�9u�ݻs���~� x᪩��*�sv������}�zV9+#Z��iLlbV|��_^�Df�h�L��!���>���QL&d�S�##Z�l9.�P@rT]Lv4$(�t�s���s����素�ÃF����(OR�j,؏�����b��̈́���&{�淊������	�]{��щ'�V�u�����`��n򰺸�,9r�@�Ë�pP:�6����z�T�"��4X\���`g7&��Z�N츪�@2=�gi��B�h�A����oB�8���̺BAB���C�������f�*�tyD�Ƀz�' E���2VW�ఙ�z��)t�}rm#�4~v�m��1LL���K�iJ�R���W����d� ��!��er�KUI�jSg����o���̀�l��+�l���]�s��15D��.�ccu�1�*&�u�#�F����Zh�p��p�XX��?�	
����uF��L�}�v�-��9E�1?���IR��<�X�����K(D�N�`h����]��������|�,�=�����y`�����S�:\z���i�U��r:P�g._��0����>�Gi���k��P��`����x��p��m����&966���~�ku"�$ֶO��Y��o�`7D������X�v��NJQUhg4"�-��g?�g].J��4��h�e[W���I�k� P���*��q68�k�l��J2�=N+N����|
�Yx`�`{g�RF�6�&�N�v�{�1�|���Ο:���1f.���������k�@ww?�����l�c/r���n��uɡ�f��$��+/����l�����)bl�_�D[P�T2���%�g(ݚ:5����l�l���eE�Ti��f��a�s*Q�q,�\��ͭmll�¹�ˍ��~�=3�F��\�,����34���u[���v�Z&��'w���!�p ���(T<9Z	����f^&X���xM�%m�	�Ev�9)���5vky LdSR(�-h�)$v�v�o�����QҩV������K/�X��a��:;��c#x��O����x��W�g��ć�vBg��'2���9��R2Ħ�L8�&z��Uv�+��s�Qz!��g
Ї��^) r��R0�<d��}�����9V%9�<O�ϲ 7%�L#���X�K����;x�E�qӐ�&h|�~N�����9� /6?���෿���lC������?�K1�r:��:��0�A���hP�l��$����g�5�I���`�YI%����g�f�΀6��4���
�f<V���U�$��\��3�b��fWi��PӖ���LdJ$�����{u+�^�M�5`!���_˰6���Ry�z1TU/9�i��P㟆��A��C�X���L�㣄LJ)���<�jU���?�4&�L���}���5i��O���I�R��3N:�&h Ԏ���Q|�����ĄH�9Qk���ǒi1�n�Ń{���؅�jD.y�\� =�~<���מ��Л�3[�V�X�71�s�_��n4���8���K�|��?�k�����s���o7��ɗ����?�ڭ��(Tf�]�H��u!ګI�t9NV�2v��R��a2���8����`w'�P|L[��8.�ɫft!U2��7��- Q2h,ߛ�7�w*?��
�t̌hTQ��$���&:�+b��0PR�e�F�F�t��,L�pyhD"ĉ�-
Y�I���4Ȃ*�UAj$��j�Ɇ��v&�R[, �O�!��W�</�h��"1b2n	(�k(&�ӏ���=�@xP��B�T��)�H4u�͗��A�6�^65v�՘T�z
sJ	���Nv%���%��L���"��S����W6�A� G��M����fA (����ރ�?��6��₣dQЄ��TL��L�zD���*�rJ�l/������P?tu:�SȔ�4�X�<���6�<.�;]�������9��)ܸ5/D!j�9���lww���W���5,�-Jx��@^�#�Zd�R8Z6�Xk�f2��+ֱ�v A<U���)���^#Ӧ%ۂ�O5�.��"7��q��:ۀX$���e�j9��~�~�2eU�%��w�� =�b2G�p�]�|�j�E��89��e��`� �V���#Qܹw_6܉�~��E��t�%	�I&�8If�J�L�P*�@��������`��0��l`?ǭ;+89�.�	���sEBb�G����@&I��*�V7����795?���H$c�A�wv��?����//"S(+]����hkwcx���<��P�j%�����E3o��w����4��0���Ϗã��wq�
��H�1q�F�跛dQ�!&UL�%�W%%<NL��;�B�RC����>��8��9�/걱u���C�JU��lZ�m:�t�^��"G<��_��ߗ5hhh ����j���ű����hWiu��@S+���'R!��&������N����9����pt\�����+�e��:eT�����4��H-�J�!b��@m��1�k��Y1>6"U�F�M}��.�t`]��N�L#��YoC�0�Ņ	,����bԈ1weq��ޖ5���abl�����������Y9�\�rA�O(A��_�>����|�ٽ8���a���d.�G�M���4�,aeeU��S���1;��W�ʄ��*������Ӟ�V�7���������OȞH���A���X�[[8<����f����z����D��W~�6^�v�f�S�����F�b\JCN�Cʸ�:��:/a�J.ЍfN�t�9X-�%<�W�+�Id������/����iS���o���\���_�I�����~�>�s/��Ͽ���O_��7���i>��4�kYpO�rrL��y<O�Z""R���	���:��~IA�W�Jq�z)�lu���[�4<�AS�g�"�����>����J,��ʦ�;���*:D�՜��� 0�`8�i�k�XYY^���G?����Ϣ�o{�������_�5�7:��D��!-� �h�ިe�7��i��}�,L,l8r�\�>	z6��(屵4�'�l`2P��D2�K����af��I�R�@� PCRy-Y��-̫�R-��M��t�&�j"��_�3~=�������&��'�NN0��R�1�p�!�+��()�sk
C+�o�j#�C�"��@��K$J�Hd��j5B�+#�"a/#�5��W�`��½}�))�z#�b���7#��Б�b�	h���dS{hSLx��G��c�A[G��r��zq?�����p�!�/�8�G6�-������>����]��J�����%C,���o~�[Ͽ��ԍ�>8�(�٤Ԇ�TZ0��)j��*�d>v���f7��&לt��Á�����pO7��;�ҕU�N�$�A��#Q1��?Y�K����`dѤ��'�����T��
<2�90ƲZ��#�:jתE1ji��'P8����<�V�ЈG��4��j�c/�Ui5�eq%bMO}�G���KI�l��h��}xģƓ�G�d����¹����j�h�8��j�05Hα!�� ��@k�3<�ޱ3v��3�(����d��u�AT�14��cJ�F������n�C��(����P�R���O� ����pT����mH�Nb���h�
Tf�����*��Z����{��U�s~O������;>a��H��**߇<rꦫ��{O�"D�F
.;�'�(dO����p� bY��-�5&<����^o���@'�{���
͸w�3o�\��ƞ���vt�hkgGڋT2����5�!���s�NWF&A6u$�Av�(Kku���@"Q���A��{2:�6]�S]�]��V=-����6�lʢ��2�R���>��XG�焇&=���F�#k�Q%R���e���S$�$�(��<t��݉�vv<�H��0r���8=Ot��;(]�|6#�k�l��0�8�c^@��LT�>��N��`_#�r��ݟ�V0=����(�Eދ8\Zt���#�D6S���6��pr�@������p{������ڲl�CC�u ���νi1 ��I銱k�n��h'\.;J�*��g�t������EѠ�|�͎S��zm��� <n��i��*T:�Zi��#�N�YfB�F�x�XH��R��6	���/�B�H</z]]��v{jvw�Ba��`����"��mCOwH~w��E����#��02:��+�zT6wP�ac�I���,�,r����"TE6)����,�۷���l��`��Q��Qa��bf3�5���t��>��5�M~�d��6�N��I&��������3$�]�d"��o����%Xh,�����嫗���Ij�ȉ4(�u�K����%�L�3*	J�N��ٳg�ibg�2�;���+~���R���ul��p��<��$�8��$���ù����k�p�ނL��>3����6���ݝ���UٹU	ӝ!Ν��X��N�'2;���Y�]�2)E'h���j��~���C$Ri�	ٟ�����p��)���T�r������9��bwAk$��!i8MU�7ʆZ�/�!���d-���Þ�cVP$�@�zI<�����������م�c$RW��K/�_��7���"����q|�K���="�?~�ۈga��`4X$����a    IDATZRu%O��Pn��Q��:J8���8j�WM�jʑH����R6�D2��Ha F�tZ�ܳ�A~S��½%�ly T��$V��"��r�(A���E�aD35�6
Z]t�bI8ZC�	0�`��k�0�,����	�N���@$����bq�U���	&L�SA�6�C&� ��DԚ��P�Y���1��	�,)�cs�QA�ߏ�P�T�ӷQ`A�#v�\��dm����Ţ�ϫ��2����hu��ڤITR2�֤�U8�k�żZ'������,����g�J5��q��ǂ��@+��F�H��S�������lw��lC:[	0�ETZp��kN�Z���S��d����R���OH镰�L�$��!Ĥ���
0<1%��,iK�u�O����'n4��&�O�B�*3Vb��(抰�m��B��z�Y�x��'>���>���(
�+�򙨖+�z�ڿ��3��׿���e�_��\P2��닏�uk�+��6wP�#�3v@s#V2��]���"�%nL��x���T���{0�����р�P�OM�iѣ·��"������x��s�����i\�q�VQ:���&~-��4��7��n��8�r�qk'��\�Sǈm�"������9S[W.����<���x�L���ӭy ,)��hn�u�`H^GR4�ݤ�E��)!���(��9�(�f0�a�[`��a'eH��I*�|����"���/�
e'`�"Ǆg�H:�CFy��İ�a�YEB`���)�5���ڸ�N�Z�����Ʀ��גG�R�$�p1G�Pݬ�9)h�	Z&�&|��� �8f¹�~ x��Hj��:� ��EV4����Hm�*a򢘾�[TF!����´ A�σޮ :N��w;
5�p��ֶ�sF��P_ �'z�2Tȥ�њ��5D�~�ά1�Sc8uz�p@�������^��^.��c�8{j>���2��0�c���������dCc�����$Y�X��d:�'e�t�f���w	��zvs^�I�����U�+7�qp,ґd�$)�q��b0���!zf�fF�Cr
�@��`6�pt����*:Bm�n��G�tEL�L�e��i,�HO��y�?smKK��j��h���x�h��"��bfn��.!��U��χё.x<6�0�2UA`.-��Q�?���S�1�`��޽��Q������D&W����`J)]��h`(�KF`4jE�ArN._���2L/�f`�3 �,�J��L���]�bY��9=mY=7���M�A��%RB��<��Yx�.��_R��VJ�#�	���Œ;;iܺ;��}�,t�u�������+ގ��Cܽ7��è�n��98Ї��Qx�N�R wqy�t&�N�QL��t�t���A��1_̉��0�83ӫX^�E�b���B�d�c2��́rD6�L���@�y�@'��Tt7�����J"�������l*���9D"��Y������gN��
{K��0��5��x�>�.-����(�2|x��et��Co�#�+�A�޽x���$ςE����8nޙ��ZZ��F��05ԁ�>?��F�U���ܻ7-��C_D� 3B����RЙ�n):�L/U���x��gE��:ꭷ�q��M�F|�ɇ04�#��\��%�[�D�h�XD�Aii�J��;wJ�&v���u|�_~,C��#>	�l6J�xyw��ti���VwW��2��P+_[�Z�0�א+�D�kF��)��w>c-��%�vu�tmue���o៿���X� ���|�._�s�}���wqp�B
�Y�l���S�Bo���$��dDSi�W�.� �� �aX�E��.#��)9���V͎u6���z��>�3��V!�2K�q�{�l���E� @���(s"��A�E��p�Iͽ��P&�=�5M`A��2I_l����8�ư���|�-�X(g6XP�jP*��@�I$�6 ��`��`q�P�^K���-�Qz�'�*�ג{�	��\ ���Ӹ���ى2Ǹ���8��������	��,n5e�M��`�i����R����ؒ+�+��O�����8�&etWh���L�O��xB��F����jB����fa�.i[�U Yij�*MG�
M�5#2���@��e�V��tV,V-\>����_����r��h2���e6�ʔ�Y�������fqbc@�$�F�
]�� ��OP��X���g��(Y�ڍ��6A�'�	9W����T�i7��ۿ�������/KA���Ǚx׾���-��o��� ��Z;�Ŋ~Ŕ�cTUd
d�V�^��B)C��:<��#x��K�d3�^^��j���Sҙ�R�+�ś-l�d��΋����k<���R(��^
�^#�d�"T���\n�t�H қi~�I�'�2�!���͹�[�A�hW$B&]�JFi��PR�S۬f١恁�o���z�H�OP�7V'SW�[d;B4�ԑL�p��/�!�X�4��Aъ�ll�ރ�(U�>�¤w����"쒙"Y����h��3w.>���F�Z�X�?L��ia6��#|d��%��.�*.t,��=Z��ʽ�(�)Y���E�QL��9�]��95i�H&��Y9'����F�K2!�?�U���=�>��Hh4X�݇�@i��YH��Іd� m��X�^�CM2hʫ���sL6�ӁP�z4��*z�lD���'�,�E�6�������e��Ƶiܼ3+��p #��ҥ65������NDR��^'��0>Jf��|=@2������.���[�h�{�G��)�ٸX`R�/��f�%D2��~���P�d�w����F��@g���*S�D����]��E��v�A�d/游7`�vU�GN�t��ЋB�mp8\r�&�5�ctr�<�شR�P�+Ι*���ܘ`����E����""��5%�xj�CC=0[U�s��>~��H�d��Չ�����ˢC����ܝ.4l��|���\.�pѯ]����	��066!�Ζ�"x0����Ⱥ����ȕI8]fE����<fVqf	�Z]�{�B��̞��l^�a�	'�idXUUϊ@XЧ3
�K� r��]����i�`5 �bC�Ca��v�N�ɋT�����N/`� �NAp��&�:�K� �?r"��H�X�	V�����uS����s88<���	Y�߇pWH>�j6!_����@�Nz{�`���ŝ;����u@o�#�m��b�<T�bAК�n��U���NL�<�p���&KeB�A��n��9-�ߢ^-"�K���9�����{[��%������c	<
�BB<���������3�X�9=)��T��x��ٙ<�?���A\�pJhO��7�w��7��/n�ǃ��0Ό�=j��	�o��ʏ�*_Doo/{�C�lg�.��q���r�7,�C��+�>�N_��sx��Y�oޘŽ�w���{/�3�G.]@�f���1��_�q�2+Lv��!T���i�
1�.���e'9#k�HN/C]��5X��M�U�ۚ��|ɖ?i�:[����f���Ke���+id�k{�?��琋��</�?��䑼��W��W"���p��E|�K�
c���s����w$!�	�0\M�M
�L�k�W�+��<��fA��D�R�F�<s��Jm�vLMM��#�J�����D�JQ�!R�������չ��y�[ ���ȕ�3��f�2� ��� ?�p	l���w(�p!vZ�N���asB��`scW.+uJRp�4ACR��f�hVS��w���ցB��t�����j��J���˺��%�N��LBbc3��Q�6?�r�\7��G;��4*��@_��ǭ�����T��]�U���P�U���-�?����De�����)�d��4���˯e�����K����R���� N��f�@>
��4n(K�Ǣ���V���T���4p8e�XFc�����u�:N��H��פ$�&J�,�|T5�vBa�I
/��l����H�Ȕ��� �l�LR�Iz8��k�J��=e�:�n�o�.���J�c����Ư��������Rw��b�����7��,_{�y�{]���&��(n5���U�-%5b"�NUN�	O}�I<���Ж��o�A9����qI��1L�� �	9�ѬϽ4���- Sw�d�ʁ�o޻���Pe�Xe<��n�mFǨ蘺ȉB.���װy�.��LFt$��<[�B��9q�2�a$�O�xt0�-H%�0M��C���]*�N��������!�旂���T6���UI�㡘A4�>c#cx��G�����ӷ���X��E�fG�F6�M~f>WF��z�a��ox��H��X�gp�41ͲA�''q �2C�(�"���LN�J�!��dC�PAls��s(���,#�%ٕ;N	�ΛW���N���(r�
��mN� �T��
�_�4`7��S���4N���A�U&&R�(�����TA+k��\_�|��%�z��L�� ��i��b�WV�NdB@�Y�f�uy��H ��ۉ�x��� ��{s������3��f�`���,�-�n�#�`l��9E�4�fH�	��G�PIL\��5�J>�]��֮�z�Lv�yy=Y�dԩ�5�<<�ΐ�m�È�]m��`���dp�bek;�8j:r��2i)d�����i�&�ɏJ9#�6�ǅr����%�-�
�}��$�=tv͸y9(��D����pphn���.�lbieSR�y�vXM���� l��5����?x��$zp��(�V��S���ū���ݽ(�/�8��gƄNA�0G�7n�����PBΝ9��.��~���+r�����ۉ+F���_�X�~,���}<�_F,���l�:	)Ԉ���@� &З��"��Ҽ2�P�s9�VS�j�Q���y�.���qj���S�mC2U��a�f��{ �Y��� .]��h��tQ(Yѓ�V�;II��\ʀ��{�����8����`g�P�=�ہ���T��ISG��[[�B3��̙s�z�������i�ǡ��`v��窮kɀ��H:�� '��~ago��[�C"]7}u?sc��%��٠�l���c�C�	u�^)I1������ya���L�:����d��M�Ш�y�����{R��V�+;b<$����qLM��u�98���f���E΂��h?���/`G�����%ܹ5/r%^��������ԍ3��N!���:dB�p��ĥsga��q���ebv�l�����u3n�\ǝ���Иff���,�2�
qY�8���*&�K
Z��
i7M=;�kZ���6�@"�h��n� Ǝ��Z���]`LZ�J�z%PN�`�Á?���"}����͟��I�s��~�#��W��u����/���������=Ї�|���˿�2����BuZ�by���� x~� O�#ͽ�Yhi�.�0;!�5M�4������#r�B�a��YeM�F��N��-�>�_S��*�o>��|)�̇�$��v��K���!��R��C�dT�13<Ou7��O�3��sf
{$���z�ܯ�6��d�d�Lɖ^�P�}A��av{$�9���D���-v�~��$��ب��OCW&�4����A>�ģ��s���K89܆����9��yhE�BI&����Y�<�wx��!�@�(s��~>-iZ�R$�BB^5u/�"9:��H�(���g�;$M�P����������	��1N�AS~��o���F��C�8��1�^��J*��K�Fy�������&�>6C��2�,^?�VN��a��E��4����
�"�"4����z�2�yʣ-�v֫y�9�t" �K&},��]+d��e+��~��_����3���(�m'=�{��?XX=����X��F�8"oR��>0� ����� a�|���Ȉ��ۭ&I~4jjx��y|�#���\�E�(��&�����;�$���n�FD��w_^ŋo, Y�f��X��&dU�� ���3j�2N���`�S�v��Q���F|sso����4��� �0٨D����Mi��?L�s{<M�K�UU���=�>���E�n�ı�����,ʮ"Z��,.�dJ�p<\�c'�f����������,��O���7�!�.ȡ���F�1el�4F�1r������+���a�@g�y��YdA ��F]�b6�Iu���)3�f'��g���7��77��Q3M�:SUȁ���EU�������*���4O��,Jy�<����SE�^������X��(%��擲�_U?K:8����l���@CmA������D#2�lI���}�j�e9D������A?B�@�\��zG̿zJOFz0:���D'��������`jb��������#�[��F��~R�/�P�0���������[ZC:W���@(��cϢ@4�5�?u͂��5�(�y�o7	���'(]���v"G��ĳbf&��׭�t�|n���]�EW؀���lH��z~a'��l|���yEOZ�瑌cmuQL�^���\���(�3�)����׶$ �{a�c9�?�B�Ӈ�H������G���プAYv+ҙ<��[��S��x�CS����ɕ�Rb��*677����d���XB�����(��q����lL�u"ɘ]ZÃ�ud�e��.��p��Tؿ$��MF����6_>H��*����+�/���z�[&T&������V"&��3�8}jn�Y��QQ;�X[߀V�Eo_;�zC�.QT���=<$!��`���ccr�)}>�ep����	�Պ��.��#IH�R���*n߾�D�.\��+�jv&��oO���]z+�6r�*$_+͵E���T֕w����N�ayL��(=5'/܌9M�1���:[,�:�x��+�ؼ ��*�X_]���"b�Q�^LL���ٳp{�R|��?�M%CVX؉���i�f����x���x����X^����:v���w���3x�ҨHV���p��}lmDe-u��t�,.=4	�C����L�v�2�7��^�( �`���O��æ�ݻ;X��A�S��n��c��/�r�gw�5�`�;��h�da �<9	1�Ƀ��hC�؀�`�É�h�*P���G��y1����1�3�q����.c2�*'�2T3hd������>�IT2G��_�)֖�ȣ������������?����>�0��̳����s��>����?��B��S�j��J6��3S��eo�c��R����Lz.�.Ŀ���Ȱ���?9�	%�V���s��"�ptY@���߷)�R�a5�c��2�R�����r�u
�J���e6�i}��V�"�IT�F��<���0"� �R�b&�[�Uv�M���{�R�E��ꆯ�%�N��\Q
�|�t�0�+%n�<��V;��(*��l����ӿ�!ԫ9�����ch�g��a�[������5%����L	sQ^������M�wZ	���g��f�Ψ�ୂ�U|��P�,�	AS/e�B��)�%���^ht����b��8.A���9=AX�~�N҈%�Ҩ�tu��ſA)�*0�B!i�nm� �w��HM"�Ĥ��f@���I��{q�Ԥ6Ve����f��j��H~n��U��=&��R9�P�I�rU&�����Y\�k0hn�Ac �*�S�]�ƹ��r��U��|?�§�����7)
�o�Y��/�����O�kz?�����F���
n��u�_T���ne����fW���Z&��߇>�8�LN	<�����Ϡ��@����fG>W���FIk�qx����HU��Y\��q@S����'��+Y� �*լ��f��T����m.b��[Hn/���L�$s�T��W���ެZ ���E`ww[:D���'p��9����pc�,!���)�4q��Ź����C;�H7�F�PW�H�fg��˯�ڵ�8؏HX���=!<�����׭RC��i,x��e�V�
    IDAT��/?���{�(�z�,>�E����8��߫"���$���Q�$����ý������$`vP:�`4j��V�H���M���\4¢�EP�Dm]uZ���+�����x�����E��VJ*�L��¹W�P��Y����P��cj�J��`��@��!�y�U�	��X�afq7n�H�����s�3��4�r�
^��[XXބ�bB�HΜ��㐢�>���Cl�n��qx���^�)�)��� �����S�F�BQk��sB��G]>5��X���!/ɪ�4d��7R�Ҁ��I.Όb�7 ��^�;{��;D"���e��̰L"#����n/���ɗ;NJ�����=�ND�.��v��H�a��?'�I!����ab|c���!W �Lo`~i�2��̂h���A��@6���̴��z���8���8��[�������\8���&�̨�d�u;;{(��2ε8���U��鱾z���M	�
�����Z��>w}���IllGp������k	�=J�t,�h�ePUM��8!(�w�(2��GF�p 8@ǿ�֫VRL�T�<F�:&~R�id��6��+S�����/6��ְ����*��y^��{��)�t�n��$Y��щ���N�`����hC8��Æ�n7�b����XY]����@�c����T6����n߾���=\�|�>�� I7����^dm��C�TCC��$�i�;6A-S��&~�heh2��d.5gƢcẠ&�����-f3�y0Ȥ���߁s�$�����ۍJ�p���R�6���c��B�ZB^�L�����R�̈�do�}����tįE@������I����&�Y���'p�t�\�[���V�ץ�nz$�ht�&���7��w����'��:fs1x\��StM6�ϯaog��cc��+b0�qp��o�ca�Z��	SM��-u�Q�n<��Vs$��̂�F�:~)M�V��]����Jb�.�1��YH�ٜ�X�6K�{�!�vNC�l��_��3HF�eB����wv��~�����3��~���7��ن_��3�·����?�%P7�l�i�.v����yI�g��N:'�ܧ4u�z�[����-��$J�̜�5�(ܣsY&�s-��in�؟��q8��Pm�!�d���M#��Z�V�S�Jp�FU�ԡ���9`�Mˬ��r�3P�}L#k]ܫ���Js�RX��#�q*rBɦ&�5*1���{`��vd+5ĳyjA9T�	����j�p��Rd�1���q�!��-��g?�I��ʋ?��?}ϟ�Ǟ�(6vvv���"�N����}�ȃ$�ѐ4m�����
}�-5-�4�̏�D���(�%� 5�2q���>��<T�at8T�*e��1��a� ��9X~t��$G v�b�a���g����C{���FƑJ�1==��u�*��G.�~�I/������٠�^G�kJ{�;���"�����ҜN�{��z�m��d�oIr7�TM��B��ϔV�
5��͢�ׅ���Ieh������g��?��խ_��໋�������ݭ��;=�'�|���:̨V���Ұ�pYU#�9�Q|�pg~�pVn�4�9�p��0��a8\حF��D�c�����AN�e���/��7��y��z���Ȗ?�5	bEH��o�C��P�1��#����*j�v�ag�6��BS�èeǊc>t���{�8e<&������l.v��~����'�4#.Jϙ-Fx\n�ص���Hw%#ЪE��21f�<`�S?733#ƥ��ff�E���މ��!؝6��A���I�P�.�����������|0y:��1����Ei��e:@������"7���*B��a��$�� }&�GY	U"��]	{Q����"�O�.��X(�_5#���,�^y�Wp��O"�m`/G���f
�lX�Q��C/AS|(T
nx���0Xc1 LA��@��r�:�ev�X݊��[�E��v;18Ѕ��0�:ݢ�7j���ӗ��<��s�w��.����܁�q;�Ql��gN�HA��W`��͕�LUa��eщD�{����\��X<���-,�1�"�+]+;2��	AC�������>դ ��G_W���"�����1)�5��ex]^<�Ky�f�C>���-0��;{G�d�^��qV].ޅJ^̪��	v@�b𤶳��v��P���"�a�|m+���M�s�<h��Po'.�GW���1v6�d���p{p��ȳ�����nJ�����p���:�)�!0h� _RYLY�6���P�9OgF�0�?{���.\<�s�{��T�cg?.~���"�\~NҘ�I�5ʪ˦���&� <�j��-�N7'kʠ�>� f�����:D����4r�����)��N��e	&K��]=�b�v�;^�u�/�.� ��%��kH$Ӣ���mw�����jT�8���
v��Y150��Pn������g����t2���6�l�����N��W�p�k0�\�5�%�\�T�5)l�T�9��@�:J��a24K! �|��`:+R��n��dB����8�b��P��0��ŹUI�&G��+�$uYc`�gE���<�)Յz�p:m�ܟY��7��U��cw[0<�g�����]�F� ���>\�r}.DYܙ���{���ȧS�h��}ｌ�	&��}��[XX� ��HP�*))��b��k+�����cd$$	�����O�bk7)�N%˚�j��Mj*��+F|�IjY�a�D�J�Sv�i�U�3R�R�IxFUo"�Pa1�t�9iU�<NX�)�5k�RY
2��2G;������������瘹uC�O�������cW����}��⏐L��ʣ��������_��9>+F�IR�'@C�C5��$5D�ǉ�'U�k9����I�⤄8L3+
I6W�L"���)��O�D�/������$�S�9��3h�y����0�_�����"%�(@	'�Ve>����J	�J�6�h`�W�
�I��4dH�1@gq@kr ����2b��3C�J�
n�.��6h-d��iDg!�B*[P
"P�;�:����,ʙ$���Fyt!4�����i<��e,.M�o��/��~��r�X[[�����G�[lu�e��>�)�uN�T\H��K�g�ł�I�jQ�Į.��J�V7�ʐ"M��.V���5����E��T̢��uz)8�5�\�:u�h
�h
�LA` lx�ؓ���X$m���� 	f��Jfd�?� �B\#��<JH�}(;eqAA͠����lh�0�X(��.�	���l�T
�<�4��~�$USh��h����f�ň*���A��"�J*V:Q9{z໿���/��_�����������k7�w>����7�{� �ۗ�d��F���Z���K�����
���V%A�ZA-�����1�O����z�|pY�0	b����Bp����*RU7t�L�-ՙ�V�pCfQP��T"�<f&��*���"[�]��Zb(��#V����V�$���F9L�R�a�������)z�=�}�{/�m.$�	�cW:¼��!O���Ȋ��th��e��+����5;x�q�dL�[oq2p$��t<�ӧ�
?z|(�=�f�7�dC�k��O��|_��+��t�- �����ŪB�4Fm��E��9�P�n+tf� ���W��Ƒ��Gvo��`,3�QˋBHRJ�#%sWכE�*��B�
��"�'M�hDI0(�`
���'����{�v����׶��(AaA�ng!�s��	>�W��lI������1:�%�DL���k��D�x�v����b/�:����
v����-��o������?zmmGR��:��ZD(CD�;;�`��rVyD6��J��-����m9�w�����/_�<�
|��N� `S2>j51�����>;e�,~�0iع�a��]����I1]E)�8���Vgg��z�A��A
���=�����B4V)]-N7G�f	¡.��9n�,���`h�W������Ww�eP�Q-��t�ҙq	m�%��N���R������E*[�YܹsK����g'a��Q"ݨ�����]�d�0��ij��p�2v�րD<��_����}<���q�ҘPe��h K�������m.���#%yɨ�KV�E���<D'���@ ��:�{�U=U7���w0�
UȂ@��}�C��@{���>tm^+��,*�(�=����]	yc�\w�ڼvx\1�%3|��?�<N\i�%�& {<nDq��[Hg2���v1C���u��+eb�Rv�I�gC+�L��R��AIc@�N��^:��r�}��Rr\TSC��[�!Upl/�f�|D�m5I ���B�ݝ835��6*U�sK2���L���Hˋ[��
F���)\�8�j1#��a:ID
���#�oB*�{Bpz��;(�7�aznV�GI�.��:0�B�\���o`anW.���+��o3`�(�������Gk���N<r�,F�0�E�P��ۋ�7��BQ�ݭ�15��:��;E���:����L�=���g�S����.^��=��`q��	C�Y��j2j6���PEСt�\U�mJ/�V֜Έ_C���K��\?[�bYc�{i�]t*���D�QD61������l����o�87-�7�Â������<+SȽ�m!F�u�KQ�ͯ=�o~�9F�H^
'g(���`��Ѧ��(�c��E�j#�R9��(W�"/b�D��Liw�#��mv��֩R��\:�t.+ZN�x��l)�E��ei25s�ҳ�6fi��/��v�����Af5�OI:bfK*���~[0,^��I�LR&l,4\�v�O�C[�����R09\�{�(q
]*Jދ�₁���Bz85�:Ӝ\�w����;��T�T M�Fh��orzb6k�g>�g��8L&�������^�gϞ����oݺ���m��FY����3OC�xj5)�ш���b�Tr
Y�����h��	`���*���M�5�o*�÷�h�b��},6;>��O����������q�<�@Y�X�Iם�kz&ut����w �T[�*8M�0U(S6$T+�\d���U�u$�Uk�˂���JQ�/Q�֔?6����ڬf���bq� B�
sQ�]0�R&�,�����K���5+�����]�xz�_��G������_�	����o���?|镟�nW�;�?��.���umE���F-IBF���Auf!�?�ۿ�ݹ�zrq#�VϪ�\������)�>QBE�.3lF�L��&��r*��f��_\ז����5{D��a�1��x�[�)j�U��Єh
Ѣ�����\d�3o�݀�܀��A%�D�z6���6㸹�R'(�+#�ʕ�Ǉ���?rUzG�QI�<8�9����s;]rCw��ho6x���C/1���[���S�&1f~���!��p�^O�H?�#����[�R����;���}F�Ͻ��~� ��:��6h�6a�k�F��HI�	J�y%���*�%ͯ��8^[G��R
Z#�P/*S�,zvKh|e�TbJ�?r@�y7����3��'�q�-�`�9����u\���LǱyp �_\�X0�`�j���jM��En��m���h,�mi�TL�����Sc��d��ູ�����*�����!�`h�v��\��{�g;��6���q���A/R�V7�<��L2'�d�M�����R�<f斱��-�`��W��I� ��"��B�o:]ƭ;��ߏK�/M�j�T�7r�d����b�I�ª�Iijt�~�,<�᰻ϰ���}��Č���@�H����E��$���삄Z1���jW��#��=�2E�X���:��lf=�V:;���a4YqtR���l��\��&�i�c���� 5�Q��:,67�&;���O?��҂L�Μm�ӤG�@a5{pp�5�<l��e��m�X�H�H�r⃠��ܙ�x���ʛ�&Wjh����[�V��`w�E�٨En�1�݁n&?[,Xߎ����eN!y�� `WQi�Q��f�(hQw\H�M��y� x�b�!��);��+{2Y����v��S���;rȠƛ�~��F� ����BowX%�k��=LOO�362���>�,fdry9<��!��bA&���0����H�[�����&re�j����H��>I9on�Lu���:��	�b�����W>����}��.�r�����`t�S�2rt,����Q�K�����	��\N���K��j�?�0���6��pȮ�Ղg�q���D�u}�oϊƟ��6�������ۘ�]��_��3�p8���?ĵ�K8��?)�4ϝ��hlNr�
�Ϭ���M�z1$��g47� ���1:��ޅ����It�t��ˉ��!Y%5���2U��|r+�6E��Z��$1�A�D3���;�U��L��v+(���Jk/��$�whI�Z�M�`�Ȃ�P���|<�Í%�|���p������/cei�*Se�R|���᳟�ut}�\�>���Ǘ���x�/�R��fq��')P/t^/���@�PC���-�ǒ�c%���B))��	�|N�T�ʪ9�?����B��N�]���ڞǱ�����=�$��e��7[��{��؆�뤃��TB*)u͚� 6�ZqU�zS�i��}�tz=�̽g���y%x���9u�4�F"��L�b�HeJ��%Y�Z�g����=3�x�g=���Y{�Y^[�d+Ӗ�I"���9�����+�{�[Mj���>2@�@}�y��>7(À��ް�����"���>�Cw�����]�[K�����0B�n9;qh����I_�t�d
ET�I��H�-▜i�%��Ev�Pg��l:�ٙ=���2�n�~�q|�����������}�oq��x�<��#�+s ��_��=�����j�C��hD[[)��c�&d��JFw�f@��8�D`m===j�ٔ�k�r@�Q��h(�xW��n'������!���ɟ����u8�����0T4�y8]ģݰ���3��@9c �����܋�����&Zn6Q�57 ҽXw��M*�1���S����a/�ͳ�m����Y �T�p:���E�� �����B&����6k����������~����+����W��/��dOO_���1���,�b$����|r����0����~~���~�c���5K%�i�����G0P��{,!���ڍ}f�aӆ��?�ƏN�"ߌ���Q�rY��@���c�ȁ��a�����$������[WP��
4�p{���Tء-+����� P����_"&b����|���7ɼr�._�(�y�:tHɡ\�QXu��u���!�s�^��'Q��H��)���b7���oL����gPT�ŅU���/�^�=]�����V1q��]HW�����8qa�fMG@I�\w�A�J�~��G�.ā��5�F��4�������^��*��*)���+�Pg,D�p7�Bt�C�Tu(�����j���u�����|��M�n�p{{.˥�����:}Лj�Llz�(��^��%	(�(��ɉQ�19:�e
-��L+lf�~E.��IG��e�(�S�X_I!����F,Ew��K���i��XҰB~�މЄ��)���e����X\�Do��hD��U�� ]�� ��
�g���.�Q�
�d��9�����ԋFE�̲5�%1�ׅɽcHp -�Q(��l[Jt����ښ�Kr|)���o<A<bCn���[�<u��|�iS��ͬ?��� ���� =�!�u~vV+eRz��r�@4֭��ͭ��؋�I��5�������p�A���~�h;76����8{���$����=Qwd��\��v�g����t(F�J!�����P��ԥ��    IDAT�".\��F�mO�!��R�p��N��x/��"�P4��߇6]��y�%����>�7�p�z�������n�Q�����@B�:��]��5_���	h=H7����x���0���"�t����,�]����I�=	�\���hWZ�N���������76>���<������`6�W�_�߿o����21�M���\����T^�\���5�?(�{img/^�Z*W�[�R6��BI��Dm
g$}��6$��m������-�ncz�B8~�(zb����`�h0ҳ����˗n ��*(��;����VtI�F�"ޟ�N^E�X��@�^��@O<~Ɔz�.u��.�XB6[U�Z<�+XODT����q����u���.�l"�S��r�V�{Y��ab�OM'�6צq���U�PW'�����㇆p`l6�O�R-�z00H�P���M�=?�KW�Q���%�E�l���:�6�bQ��P�,��~mI'��kͷJ������4���D)���	�R�=���4[o��A��C&���D��k@ju��ۿƭ��$���@����>����S�
f
5��ӧ_�_��gq��s�g�j��?�#[�9@51���ӯ^�F�Y0nx=!8�zx=k�eS(��p;�yD>�D)G�a�M9�0|��/�xw�xH��NjG��V��p�u"C<�M�ep 0�mY�*K��5Qg�N3��;TY��KW��q
Zmpz,�<�����p�-!�K���M�+���Ľ>���I�g�VS�ź�Ʊ�/!O��liR/�_(jʦ�4�-�u�v��g��:�*�Z�
gQ���N:$ϧ�߉�H��;�����u�z��n��FrE� 0�.��]2q��?Ӱ�ׇ[ѣ�F(̾G���:��c�<��ZjB�s���N�YI���ӫ�t��[itw�*M�ߛ!^��G���-
-���/��7�'Aq�Ep��>����S2��I��h@�ٱ�5��"����6�/���rڊ��6��xݰ3 ��b���\����׭j���<lt2�h�������j7�-�?�R�t�+���^D�T�%��-"�8�����~�����#����ۉ��w_�ݓg�}4�ɹ����3��r��j�;����so}�ņ�s( ���ƈ��(A>�����"�nk����X n� ��SV\Tx'I��5���
���� Z��d1�wqXmco]����
[ȯ�!�x($a�Kh�v��n�艛޴�p;=j��V�<ٿ��;��w>�ׅK������Z��cPR�|x#�^���������؁��~�����K�p Nוjx�W�rF�	��8�Ο��WO����Ao�~7: /���E\�v��O��}蛸���Ó7��mC�]B�~�Ssj���"y��j� �c)9ֈ�-�63�,. u�l�lV����a���S\��	���|���6�<�_��]�6P����y�)<��7!g�!�͊�D�r��/�B���ؒrD.)� ��Jt'��g�I�#��g���vV����ml�A@M�{��04@���
A��8��kH��R��\6�Ю�+)Ģ]x�{e��r�ĉ$�u���8}YN�����\w�=6�2�P�L�е���L��Z��m��l�X<���@���R���n����`&�	�(W�*�m!�����u�9m����QD�^=N�5�SM���a#��p<w���,�FI����z�܏ѱnafܪ���q��YT�y����	!J&(Ё��y!���iTh+�h*h�.8{G���A��Ѵv�D�I�KXXY�{�ky��c�^�R�v&�����ߞ��h˥4�JQ��{��&���ifLcn�&�8�#�� ��(��6��/\��&R��&�~����]�`l8:��X ^���ڦ(k�&7mD�88��@"��ݦ��
7�:�E�C�({���#�t�J�����R����좾�'�]wLbl�K�[��qkx����57��sh�t|o�b��ƍ��?����`/|�ׅJM6��bYu��rR�(��V���N�+�8sᒆg��#kD�	��^7�����9���Ǡ�M8�}�( �C�G^v�HP(�����B�s��eKG��h��aC<����7�Z9'�ǥ�^>u��,Bј�Rz{|x��{d{��2�n3�I���&pp�}GН��h�G����~�����8q��R55�>r��4+�ƾ=���f��@6_�����+�p��RQ�ۣ�1<tl{GGD�=w~�n�"����qƵ9d��/�����Q�Y�CWo�¦2�i]{�]�:r[G�]&g"���*"��d�ßلh�����lmwàJL-��͹뺢���E�JE؈�g����~�7V��/�=��\T�
C��N�t5�7?������p�t��E���N�:%k�;����<���142 ���8�?���*�Z8և��q���{��Z���2�����H�,"u{�lA9�x�ۅp,����OC�D4���i�1�v�q��9log:�u�Ă@��l���['|S��5���1PM&��^����SO=���_�<i�D�S���[��d�'��"��I�TZH���hkR�<��3y��I0���d_.MEΖ�\Hsd6C��A��C��f�k�Wݸ�h�_{�웟�G?�~�<_�.�/��g�x��������S�>���
��2��5�Ͱǃ�VRtY�����l�	<��F#бk&�N��i�܀�Ռ������+{ፔ(�|��x�;ގ������(�����_����m��A�҄V��-���]0i��9U=j��J���zE�0Jcv0@���4��yP��
��N0�du�ef�D6��>�'�����A��:�c2���Z>B�(�A�h���L!�\m$���?��w����ѷ�z�����տ:���ݟ��������~_0���^��P�Յ��ho�y�3x�[ߊ��<ʥF{�34�[b~��A���YY@F���"���6��j�M�n46rm|�{W��Ssȷ�+b<��v8I͇�^v!GN���R�b���毢���yX�,*�-�]o:/��^x=Ax��b3�z��F������W��.������ܹӸ>u�}�Eww�^ ���B�7����`�_�V�D�U�hH������իZ�ix�<��x7���pkj���?��Y5j��l�(�V�ڠ���=�$���u�����ZB�ݥ<��(T��:�$�2�:�����gs�wB1����-dgo�4��'h#�iӋP�5�����ɼ4S�[��p��K��Z�jjM����	<��gPt:���%j���Bn�\��\�́&��d�H�Մ�n���X+��;��{F����P��v*-n;�L���\�� �ph�]�t����+��p�ޯ�(!��]kqa�J[[fM0/� 	��:y���XD�����h7Q,1�����&p�=��XH��{����I��N~���r���N�6E�iS̀02���016��_"��o&Ӣ���Cg��^L�	]��ɛB���������v�K���*�\���r~ G�2��E��Kl��Q��\A���P\K�\݆��\�2�d�M�.?��
�a�L���䰐5�p!�����<���P,�g���{]	�~Ձ|���[K8u���Q(�ĩ����kҨ������w߁@4�r��d&���.�Q���D�;(�Â�$/,mjېɖ��e���p/&�a��K�Ϭ��fM�0��6�
��"Q�<�MLGk+WsИ3��sT��)z�|x��1�X�*ĭT�a�����2f����w�ȁq�����VW�nh����`?�;&��k��k׮��;44�=�#���_"E͉��$�g�4X����O���E�C���\�����*����,��x=��l���a���(A�]-E�&��&�Z��RgF�grb}�~���\˫�������sX^I*o��s��6-�����Ǿ�.�v�)!R���s7q��e�*5x��(9ǎ����	Y^�v���D&߀�t"r�ر}���xS��6�?�M���2^�x�iz��Ն�����D?17��6SILݜ�����̰�zƼ��}�=pH|����8��}�^���~PGK��ӧ/�,Lgk�хb]�����o�>L:�H����5�t��u6D�e��GOY�h[�7�͗��\ǎS����ȟ��}�@�Mn��Gi'���^|�����<���/b��%8��/�@_[����!��η�矇?D;�Y�ɟ�	~�������?�>��_���Q��n�Z�����g�.�A��o\9�pH��bn����]j�m��`�5�T,�dO��:�Gy;I����P�?�0ڰv{s��k�JPH�&�,�x�S�L�A�����Q�t�����=�U�E�Y�a��c���G�'#�/_�j��m��!��.4�����t#۰�n��nwJT�PZ�6ɴ���G�ڒ�5tol�2�<j|�D�#틉��D���t�6�Q��7=�$>�������ʑK�ۋK���?���T?X�
�|����@�S��}�����\��w��x4���th2!��\��	��>��-���\��Z{�!��B.'-��������'?�w?�<X�����������7EO�f��zZ�2�M��S:!�d3�yM��h�2�/��75[.[�R᠖�XLS�
 ԕ@��B��_�h�n Q�>ޓJ.�6�Zj��/t,�5P��-3��3�nn\<H���khW����﻿�k��O��{���&��������7������@0��L$�?��֜��pW��g��'��۟|�z�s�_\���&�Gp��a�u��Z;#���z��XX\Ǟ=c���?���(�U�w]�RT��@��.e�����ʋY~�mx�6��<R~oa��e���^����V9P��K*Y�[y
����^*��Z��h?���7�]Ͽ{���t��[��IhP�8��2׋\I���,��~m@�"�jŗ��DpY r��Iѫ�hc`hccc��@ţ	�ܚ����7���¼�
l@�^�������4��w?|/�V*�·N��g�a����MN���E�T�aw����đʲ����ԗ��6���;s0��!����1��ա!���S��2�����������X�������oG+��JjC�aD��
x��o��ͯ��dK��v��.8h2�Hģrja�o�Q�����P�\���RPdY������~L��cRu�v��Ҿ�nT�%%�nl$e�7<8"�(����ؠ�)lm�!vhg"l��r%��D��H ��N�̙��Je	3�,&t����äu�N��6��Riz���CW<��Z�Q,ױ��.�I����p7��5a=�X������ȭGE:B�7 t}'�|�".\�!k־ބ��D����f�3���P.�������˘����Ӌ��=7��d�����w�]G'	�P��D�)�m��1���i-80��ѻ@vO>[�փn_3k8u�2R&�a&~R�W���n���{�����
6w�q��i�����O`�Đ�*��PJ&�
e�������]�����@�V�m|�(�73�xe�Ԏjt!/U�v6]~C�ik � K.2��N/�K��6�{BxӓiPͥ�u��Mk�n-�)C����"%l@��?e�5��|^sn�Ƨփ����k�%�<t��z��c�kۆZӆ��g�깋������탃	Nw;������]���ƫ�a5Y�7�v�RW�E�|)6�y��)�d6`�-D��%&Ո��ha�� &'��u��3��&c ���v3s���Y֦�nN2ܾ�t��<��1���fn��{y��2^=Y��dDp`��;*�Kn�+��}4��s ��7V{z��V��}�(?�����X�d _\�U.���Pw݋����S]o)���kHgKJ&hsםq�~�cy9���^���SBF�x�A<����������n�7��G�f6P�z	��_6������m�� /�x3s˰��p�ʭ'���-V�"�1�P:5�u~)�6μ�fKN
z�b~��B��M���|�]<�/��H�^��IAk)����P��:�_��G��U�ş�ٟ��?�#!|��ǯ~���~��k�26�r���	/~�%Tm����vp�J����KX-��$����P�g���D���l�#��H�v�{��rH��n����0uc��9�&QS�|n
����b�/�лH����(<�����٨�I�^���>�F��^n��dm���k�1���b���
���|�י�K�%iA6�M5��;B�I�蔛S����Ԩ��a(�5�<S��|k��crRx�r`A9�GhC��c� �w�-�Z��~�3�5�I�H%�3���T��D��h�X$�I{�.^�$@����PD�����M��O���_��t#�B�p���{��f�.�S�}7������m�|b�.��vL/��_�&~��SXZ�D�}˭?�	k��Zٸ0��h�`��M�=.�!�w�V��#
�V����:+D�����9Q�h=����8�N�ϫr�l���%��u�y�#���C5��)�7�46�Q¤3W�p�K�{z��[{��|��~94�|}�������ϗ�_���s���Ð�A�B9��c-�ް�>� ~��?�W�^����/�;2��{�|�7�����O����>�����������E���� ��5|���8yqC���=�i�t 
}5�ٍs�,N�9�=��(��}��먬ހ��Gu�▬_[�찹�j@�~��U
"����{�������O`gg?��06>���Gt6n�|N8-��3������Ŀ+��^�^ �TQ���lY8%����!�����ҩ4���q��9|���b.J���O�'�A�$�Q�\���N�s�x	k�.�{���օ7��N�p�!:T�+�9��:��!x�v�N/`��Z+K@qG�͢����5�֘�M9-[9�Q�-� �/�u$OOA3t$!oN�̎�!ҷ�����|V<�ō5����+\RČ�`�1a �ܸ!��(�#�1;-��=T���
��F�������<D1�~P��`h�mn(l�l�ȑ���R��O�6�� J��g�nd�FjQ�Z͎<�|���l�K�*z���g|X�f~n�+�2�pr �������^bA�1ͻ�&�⽠�'���~kb}3%�W�}]���&%&�!pq뎭�,�;;�Ts(FcHm�p��nͮ�VnH((B_�ī�A��)�u:k���@*����T2'�aҭ�m��j������8��<�yn��ҷf�1?�l�e{�q�Gd2���B�L{6kIܘ_B�L�W<����k�qdr?x�.���L�.gs�t�2�o,���w�}�N� A��I�W߬��'��沐)��āz����&�N�B�ڔ�;�	��ٴ�������19`;i���6Y�\�Ku�����D̃g�z�J��D�k�SXg@��2�9���`=�߅��9����q
�(kv7�����Ü��H8,������Lm�_J������_D>W���E7�٤\u�q��~�\7D�:{�f���D�X�p'���*�k��.��	�i8���9!{F�!��L'ക��9��r�)s�BJG�L�J�\I��멌�ݑ�c8zpng�4;f���p���^���������q��*^���r��e�h��`�������`����N.�l.�ͭ"V6Iwh#��"�����0��1�B��������qk�$l�`dϸ�����P��\�0���f��=��]xӳ�Kߔ��P�83�����dJ�,�v}ttPg����> [�Sy|�;�E:O�"�' ԕT<T��N���_�!|�#�7���t��U�P+6�-_�9[u���H_�:?�.�P    IDAT�~�#�76ej�ڴQ�U���ˢ;�#�<�g��D��_��N��7��c�>�}�=��Σ��R$ˀ��|�+���� W�����"9�y�lΫ%X�"��n����@,��XK�Bf֐��?�-1�E��?��t)}�v�?��+�|���!|���[&g��iOO=�1L�&ȗLn��3N�&߽ 7�?{�(b���a��^�{�|�ZI&����5,�na5U��V�%�[z��E`s�d+J��~���-�<�e��U)�Z,�U��Pŀl���{�8��'PoYE%���k�{�������@?��cʃz�嗱���A������ ����+!��\٫���3�"��C�B�����ζ�����{ �9�ŵ9d��s�m����0�N�����{	�T����Q��M�������~.��Z�K�� ��'~_�v�rڌ����M� '��~��sΨ�`��1����w%��Q�9˞�Xg����v����&��,�쌈��hol���S�e��q��l�A���;4�����ǟ8���Oz�+�Ք��~��O?��?z�ܕ\ސ�VZ�@�~0�]����COЋ���>�� *@տ�J���o}��x�0�������A_���p��p��x��''�w| --Q������' �/n��������(��
6�Ä�-�_�QQ�Z*b�L
��%dWn������7����{M7�+�B@�@�Y�K=D_c�x��o��� nޜ�ɓ/��s�G�r�of�r��-��CDkWX���O���k�1�#��ѿ�_��X?_�~�J��J�"�J�TË/��s�"_��f���O��h�9'�����?��|��QĆ���l"_k��l�ؐ�J�9�"����F��s+ظ1���2��-�*+��V��N�!g�#t�Φ�H%1��i�q���y�f�4}7���A�P w��a<���camղ��w�]hR��N�b���t jp�3��۩5;?!��Y�YX+�l�x��/�W �Qiuh����9)��=�Ji�AW�0���G��N�99����۝ύ��#6�M��ɳ�|n���ķ��Owcmø�8HW�n�m/y�y�$���T�X��m�����T�O�K_�RB|n;"A����GW��Z`}3�`�I�Do�n�w�PfwL��{���A�E8O�9mE�����N��n�l��8��*s�k7@,va�hFG�b�U�-�a3�#q&��:��#�\,�P��!���,R�Z��PKK�fn{�\ݱ &�C�p/�^���u����tQ�؃���`�ǏZHn$�2��	:���ΡTm!Shcfvs�B�v��T���f�%����5��g���/��yy�7Pi	���7܏��4f "^���6ֶ0���,��x��.�w�9a�B\���Ϲ\�$��cBї�VD%��E_O����ו�5�6s+��O�U��'t�Ir��8zd{����iy���
N�� ���I��W������U����ԁ�Y�W�Dw��Z\`�/�Ѿ(|�|�:~���z�&��e�ݩՑک��Ԝt&L�C���@r �-be}S�}���XDMb�X���4�M-cn!�'�:T-��t�1����H\I$�@�ʤ94P(���,c3��Q.�16ڇ����� ����k?��|Y����<^�~�����H%�8�A{fA�Ñ�{��wb�/�v��3l�%��L)l%71�w ��A$����b6]h�C+vB[mz������������^�~q P#$Ӹ�N�"U��tQa��6\6x)O��U�A�e���V��$%�D�}��5����б����8{�6Rk�;m:S�{�q����'h�������X�)#W���ۣz�-@){��������E^x������ɟ�~=;pW�y=礪�]N�/�!�������'����z�!b�������8�������	�	�\gϞũ������-���	��|�'q �=����VV��h8B���f�qaj	s�i���Pk�`�D��Ѧp��[u9�1혯+���ʨ�*�*��l�tg�Mܜ��$�M1�N���`�z�(=[,D"���BKE��V�Q�0ŭ��	g�Z��Β�yRd:[�g����3̲�\)/�^_o�1���q7�(^�p8�^h��TAn��K�����{�g���<nL�Ȍc+�G����P H@0uY�fLf�AӃ]g8�ln8@���;$X"�إW�5��Q��>?�pm�Dj+J}���Ѱ��.�(X�"���V:g�t� (�Nֈ慓�W'��t36Ԭ�Ԩ��@��Z~�v߱����������_����n���/|�o-��c��d`��/��Zi�Ǉ�Y�#��ޣ��wcs��p���#n��Μ�o����X�����z�.����<��#����p����i� �ZХd_��Y���*��n8�	�0��B����b� 	&ZLgm���+�H�L���r+l��m��2��Ku2vs��f1?�ч�Ǒ�	8�L����'���k�q��K����x"/&Zh��vP\���*��(�]z������HS_���T��y�'�I5���I��H��f��r�h<y�Q\�>����{�ɦ�q���p� �==�)�-�_�G���M�M<��}�"�/#S��4W��K�G��`$�&���/>��W7�5;���2��-�m�Z���&���6=��QR�)�����2�0q]�F���rb0�	�Pg�ឧÓ�y;	��꒸�D�����kȤ���7 �NY�����e&]r�jԘ�Lv���:$���*�3��5�mU��&Փ��27Pe�!��i�h�}�+�+B����f����B�m��h��fɤ7�Yc�E�^C�0(L�"B���{��w2��K*�����s�"b��˴a�
�;�؝�)>�a]�f�J����I�Z*k������N�|m��R�����l^x�bQ���N_k�ܓ2���%�{/+�O�t�X[W"�%���VY��@~���ִUQH�eC$D�}��Hܶ(`��@��NrD�����?��3���>��w#�P.`c}���L^V�]]a�yd��p���mm�=	��.�U���!��"��bqy�TҸ�9��QP��]~��zw S�C��C�`[ݴʅJ�z.w����c���u%_�b�v�k�_e-`C��_"��`o�6W<p�g�`�;@ʗ������"������ � ��RS�76��-�<������{�g�^0ɕ����^�����L��L�zG�ʍ�|� m:�d�!1���u�h%���WNS�X���k����-T+�a�h��F�	:_z�R��05���W��;�G|~��B0��V����Ts���(�������XZނ�lؙ��B$�ơ�Q%io%ױ���p,��#����2�V2��Ӯbh0��;�����Ŭ���V)�-V��GW'�~+�*��(�׷e��͕�pǢA��q��^nx膢���d��P*d�z�?��&7Wlcfq	/�zk�����YM^$nI��A�U+L���^@�䡓�{�瘎F��t�0��(�שp��D��[W�\Y@3�S" ���ZNju{meh}#[IwЍ�l�>��;�	���[�/�L��KI̯�1�̠��A�%�	�c�!�Q�P,���~7Z]
S������.T[����%`ǆSvʤ���X[��O^:���$R[e%�a�888�'�x��{16ҫ��g7��O��������kS=�ΒU�-��t����)���b1��w�_Amd@\���W�^���6R��V N?7~��qC@�n�^4�#��X.)GÀ�&Ԋ��ͧ��x���W ��B�\@�L�h�AQ4s�8��>F�s�r�KL屔�:�Xw	n�� ݔ���q���S_@=j$y��O���h��۲�m�ͽ�����{�s�����uN.��,����$���A�Dp�l	���8f��+�~��-cC�m���͊��#~?n�M�Bj?�՘���b+�G���9�"���S�РYs����F)���Ђ_�
Y;�?6Nf`� ��ِ���/��6-�
ET2��C���o|�O�_���O_��W���5Xo׻��g�K�#U	:)<��S+�=$�E�O��L|:���O�~���r�ȇ>�'yS�oaui�Lbt0{�U�D;�h;�Yv���/�<~zzt���2�l@-�%�DN����*��א���Vf	�m�MXm���̖��' G#>� ��x�s����8vҫ�3>"����D��M]�׾�Uy�9���;1�a��������ߟ(FMr'��}�eH�c�U*�c����N�}}��Ў�bjH-��7�
�a�����(,�c
���pvs6���/?�o�'�5B�s�m;�ng�HWj���E[�5�ǡu'����J��mV�к��Zf6aw��p�Ԩ��Lb&m�F˳zYu�8u0�e��v��@ECA0m4�.�=���7��?�fЇ��E�km]gڟq+�3D�h1���A�P� �P���
��z5i 5�4�D�,"W�7u�(oVԼl'R�;ऋQ3��L�r�0vkL�&�����!�=!!��@���^�;L��u��7�PI��������Xx�/�ntDO���x������Y`��	#� [6knԊt/�y^t<�Ӽfk�B��b��Yr��,,�m-x�Ɖ�F��dRAd3h�/�b��1;E]����I)����
lV���j�x ���j�!���7:�4��*��pR�h)�k���.^�L��h��9��rsXmT�`F�hT((��I������R~��	$m�jHe��U���o��g�a"����^�,��?@���il`�3gǕ'[$Ռs�]�t�^�5�M��t	�2��|��۸uh��q�Н�I���8^�
��
E,.�J�GKaZ?�U�@!���t���9��g��0R�:����׭!����R	3���d��8�#��46����wŨS�� ��z��f�)�}4�qYmD��7.�N4h l�j��d���^9berUl�1���7gQ�T0�Ӆ�xD�!��EC�̌�G5�)�Rm`}-�3� �� ��{�G����@G3�!��X\Z���w�aye7o-K�K�[6<3Ba�R��"��J�&��Z_�6`��c�#�S��joI�ᯧ�U����	�Æ�ϩ�� 7w1�D�1Zs��/���o~�P���,.ߘ���m��L5i��wM�(Չ7��-{�1)�ry3����x=�X���T����DnZ�
An��X�v	s���/NnS�dicy�Y�Y��J7`sS�܂3��k��12:��DP�(u�z=���w�+���:���u�`�I�mV��0��`�w��z6��!��DTr�piyl��E�k�PN�Oבc��^>qFt=f�x`�!2}��A|���3oz� �qF�ŕ-����>�������@( F`��Rt�����YR������?D_����n��秮azn�\[��nf,9�ږ)j�Q���&��5��� ��9�4�S�M�#Kpi��S�)q��B�ZJ��'�8c*ěgX�[���5
�,��JTB�͎���Iu�؋s3���@q�<P���6z@1wx��}���P:�W��������69�8q��/`C�n#������G�7�u{F��j�ag�Hg
�����c�����6C�J%̜7�c��GgY�X����v���r���I&��E��Yd��h�+^v�5��$UAz�I{�7��a�w�������+���/|��G-����W��_M�ι��������~�W�w��n�o�^�ỳʜ%�;�x���]^v��t��o��G�_������~O=�4nL�b��6NNb�;[���@��U��߹���ZD��M�V�+���_n���e��ن�U����M�G+�4v�ZR��@&I�;r��FF�����h?y�>L�F��#[C��BA�|��������:no�i���C18:�r�,J׊���6��BO�KBTL�4��|�on`ff���G#r�����Ӳ�V�b>؁W�| �+'\4�,.n�o?�u|�K�Az�Gl��߈�G�V��T���ݍ��|`U
�k�E䆺6���D���$��MԶn��(���3���ǀ�z����(p�Yxz:I	�ߓNmrR���łU�6`�r�q��O�M�{���Kj���*$�ݮ��:t8���jX�x�4J~
�ZfJo�a�:a��zE���T�wRW):֦�n8���w 
�$&b��v��Y*�B�<Gn�ZlX��_ϯ1V��Y� �˦IJT�,�\%����n�D���i�P��q�s�p�<�mt�J��˫À�{�R�B��1"͖�x�~"k~Q��BA��D�ZE��EU���ϯ?�AhDZ,�lɝwj-��dLׇ��||�E찷̪���(7Eh�ժ6JmiF*rKQ��2�U�&Y|�����d3p���U�X�א����9�M蹩7�`��磍6�U�Ɖɢ
b���B�I+MRY�;F�BX[Ru2.#v}f�C3�Q�F6\^xv�5�+n	��:A�tk7��V��&��IT,Qd���EUj�$(G#���k[���g2�|�����E�g���68�"��=B���m�'��"ڤ�x��0Pò�X*#S�+���ݯx�����g���>_r�0����lH���)��C� 72lH����E_ODw���9%�,�+�ftd�bA�ӵ�4�r�g�Ъ6v��w:���qە	����i�8ئ6�)�{�G��`����{G0������Ï�+N��˳�zm�2�E]�=��0�߭3�i��'��z��L+�:�-c'K�Y~L�|��1u�T���,lm�ò�q��9=�Px�.�B��ظ�?���+k�q��y�n�����%��ѥ��m�I�@��n�#�Ƥ��>t�a:b��|�)&	�`��
8�5�x��Ν�;��Ӏ��7�1�m��`  ����S��q�ȱ�8txJ�4�\:���)T
ED���=�,\�\]X����W/WЮVp�1��a�`�LsE�^���U�M}n���qQg]f�m8���VB<]�fn-�qS�N
A$����}�}����0عn++I���~���3��,SK��r�Y��J��ݥA���
��Ό%�ު#�#�7�`�S�p��"6�*h�T9����J�(�kT`�Ƴ��@@���&6��"\kw[�K��x��1�e.�Z� z7��|F��`4�Dw���*�T8�*W�j-Ke�:f[��,tB֜���'f�o��tHst�	x1\Qr+�\���_˚Đ9�6�����i��H�����nMϨO(�j:�<W�uB�.�N�S[{��U�F[���Z���?\.c-4k��94���n4}n�A�xF�W��@A�E�#Чs#���B՝�(��A��5���P�v�&)I��<�t�&��I�|��W�#���/e�'.�|�o����|�g<L��p���8����jՄ�G���n�B�mo;_�7���?�c����C��qu���i$p�V�*��:���\������������R#���:Ƥ`6z��rp�ۤB��]Ϣ�8�����,�4PM�Ɣe��J��zʂ/�������h&XN�+@"���ذ�9ZԘ��B�V��3����-{������w��p�\&��Ԗ�2�A��.ٌ���t��/vv~���oZ�q���׃�?���, B�Y(,�q�^G,�%���SW���w��]�71�����0z�>4=>��
�9ikW����r�hK(JS"���ml/o������;��rp8���e�UF��`%6Z�]�+1�D��v�In��ņ���@�oN�    IDATR�u\�����O����U��V�^��X�a�6C��΀ m��5:v��\c���47h�b
��vJ�m��,�?iPoٴyb�Cx��q͆��(A6�w]�,�a�,0��D:X4i5� �&'jU����f��@���RY�H�O��]h6�,~-	vW��E�r�,Sϻ�&�M��	�H�`�%�+�6�w�:Xi�tآUi�	.�W�|�=����A�)Ho6��v������q��z�Ɔ���_�o3)Sl}y��_�kb��af�6��č2�hK4�b�(zj� ��ф4p���U� ��\�;N�����ψ~�lN��+�h�b[K���7��9�0>��$��g6E�I�5��y�8-�I�$����8#��jD���2[Z���9��1��ְ#_����`�*]��6�k~��j�"��y����J���߯AA�.^�z�r�FQ�:��k[B~���/��CJ�.��&�6��6\�rx�@/ݐ�@��L�(��,j`0��Kg�B'�f�Ϻ�h��,"n��+W�re�}�AN�0W��2G���I�i�Yu�ٲc��F	M[	� i	�*^W�[��H��ȃ�r��kܠJ٬��^ZT�]B\�Ɔ�����i�}f��*e��Dġ�TEh�=�FW�p@�n�]���3�Ц6H���a�͵����ŜU*EZϖ06�/KUr���5_*cyeM��`0�B����-QR}�(jM��tt9"4BJ�?��[t|k�Ɓ��4�Kb�=B"S?w������^�J��x �w!����ԙ�@>/�e��h���.p�X��y��Y��|	tE��±{���� f����+/!���&�{	������p�GaE�J_�Vr�Cɀў�����u�^-��M	�%�,�I{G�x���n��G�lD�NRR"qm����(t�����E+8��4Eܿ���xX�#�(u��yQ����e���Е� !�;�@w"����d��>o��eYX.�Q��r���2.^���z嚅Z�^�BżhUT���0�̨)����;�x��kYq��ɦwMzM��Z	�JNR>I����ހɭ��p�Qk��=_(�J��f�<9 Q3�k�� YI��@�10YC�� �`.Z咝`��8|�Yb�	�n�
#t!�Q+���>,����ի�5=��	5n�&ưg�z�����2����|�-��Ѩ�����9�,�bs#���pL�'�I!�K�������I!��+}K��\�Z�rkM+�LN4qY�����@�{���I}g�䃽2|���r���C���'?�§?�˲!���_��/��_ͯ�?�?8lѕ���۱/�zȡ�+���cx��C��B�[Z���*��l�~z�,��?�S��?��O��c���)�5;t�]A��"4;�O�����VK�KgVQi�����s%�̓�֌D�y�y��'GGyե)l/]E)���@cۼ`z�8���n���HK����(�M��݇���#�:�m�%똎�sy�ng��J [�cemU4��|@Hav+�l6��%c,���(F��L�YJ�_1��٣Mە���r8�������G��*d%�Nb;��\� �Q(����:C�pq���?­���6Z�.Dz&1|�.��F���A�I'��u;�,n�ӹ��i�Ë+(������vnNg��[;�&�R�J����+�5��e'�������@@��r:�4�_��Yi��v��7�Q��ߍ�n$���(��Η�����w�9;�������p��i�,6�l�L,<z����T��9lwH�����P�<'0��;�|��L�RV�����F�5n*�>��#��a�T"ϝ�ݳ�Z�mZP� 0a)v��4��#����y����s��i
���KFg��aT������)%�2���69��Lm�W��;3��C���c܍Z���^��\�:\(�gl�+Q��ܶ���v��0�9D�% o�X��ckɖ�{.r�98)U8r�^�wD�uNK�q	��y�F�+or0�t""����Cz�^��8n$v7�&
Ղ]�L9�^8�GVj@sD"9ᯅ������n�L�5�	>����Qd�U}�X�h�D�Q���jǃ�8z�i����i�E����Aت1���F����6�L(U�h�׀8�k�v�DU"tD��.�Lf������!��T�����i.h��-�L���b#O��ZGp'���B��wJ�rMJ����RQXg#��;ͦ�N�\A����I^�C�W|>�D��"l�ꨁH?��冻懣�N�[�
�<l�<��d��MA���5]A�Z�;��p�PPXS�i	@"�c|���G�+17�(s�9:�>�cQXn�l�BNg�*��|n���Fw�����~:ƴ�(3���.�W�	n�8�r ��tP�YRs��W�oz� }/��~ؤ����`��j0�`&]�Z�Ӌ��d,�Mo�g��)�&����]�E�݆|����u!l51w�4��x	(� Q["���$���fsh�"táMu�X��½���K?Ņ�'P�fD��6���#�w=�f�>���ܼ�����(�6`k�4��}��v�zI!�����t2t
6T:��1Cg�H�����a�<�[Z����7�E���+�r��tI"@H�>��~�Em���VC������E�s��7���t?��X��;�v=����CQ�\\�Y���%$Se�Y\���H�0�A:�`eB�����hvx��~����ؖ�٨���F����'�}n����;�2;Y��e=[Dwӛ�ً%Rx���
[噳���-�V-,ҬS�8MQ3@ ����%7�d��`�N��|�]G"��A��:�[:@s�z%+�w�O�晠IoL`h�^�&f�N0��?��giӀ?lU��Nnca~Y���7�07=��[2�������`�Chv��̷H;�@��%�������ZC��� ���L�xS�����Td�m�8��̽g���y%xnΡo�΍ht@H0���D���9G�ؖgj�ry\�k��;ikf]����lY�i�G�hF�#� � rjt�����9�m��;��V�j6�����{��9�	�2j�d��[<�k_���<rl�b�f��>��)C��3��|�������ڱp$*����J+�K��ܔP�gob������qݾ}x�ݷ���/`[G7|�!̬n�����j���o���	�?�r���{���+��c�&jؽ�՚�8�X�l��ϝ��-����2H,dNX$�+�� ό���ud�Ϣ�:�Rq�n��q#*���6�p����O�����"8�o��~�����X�����1]H��{�SW���+.u<�5=�龲��.4�e'��Uc��Ӈ���h����i\�tQZ��;��*t��9�Ri�~�x�z�߉���}�ML�N"S̊c�k�^<�������W��o�E��ĥ�KX�,!�1�����ߵ�k�(�ߪx=�q�[����@HՈ�>�l`sa��e���&,����$,��UψSh�R>��J��`���=6���@r��rya�WW�}x�{�|�����X�o��&��(7�&Y�֌�X4��Z	"")A#_K�9Ц�0�Bn��)�6Qxn׽�W��xb1H�2qyh�M1�l�m�m�cG�Ĥ$��
U��;�∖�S����l,�b�V5�r�)��x(�v���f��87>6tq�:+�*pX���0�rG�|E;�����؜J��J�H�66�!�ֆ�x�bE�8���Q�16.��5ΐlp�FWA6�U���S�*Ő&�Z��ɻ�5�V��4���I&�B�⪐k�l��+��C���cA1_����k
����Lq�]�ʰ"���9��ōfQZe��|�|��4�D�����M�fe��{b���#�J��)p����4��9-�$�<� �r���Q4Ά�19��,���GĶA��F�<p�^,,�h�(��E��P���C�p$9�ֺq�b�J��/
�Y#D�X��.D�����x��a�q*Ģ��$w�礞�^m��5o�ې�GGV���kMp��L"nP��\]iz�~�F��Ԙ[�=��$o�M�"�(UI[(	$��E$��[�X�z�� m�-��)C�fe6b>�*����bC��Z��dl.7Cԣ ܸR��v
U�VXS�h�\B8ȵP�0�^�l���2���,=�� ʍ�l8e].	�6�pX�
	��z�t:��FgG��0&���_M����F�*�IM��z��*~;<ހ��,n�a���L��Y9l��ɹ��do�Ci-���rq�ܱZ��,,	>8��ٴԄ�G�V̜=�so��3z=.(t?�>b�WDL+�ȷTaWnM��7�~3��u�&/<�4N���N'�.�4Y�D
��N�v��=p�V�	�ؒ�@1{���ӂ�� ��|��SSF͍&t|f��Z�j���	(�<Mg����z�݃ٹ%����H&�؈�P*Uu-���L�m�N�āa��t
����X,Bw��=B>�@�R�Bf5J�bIgd0���:gE�w���cf~//bc#�l�*Z9�Y�jY�4e;j �9w��Z�
�d����9H@��ԞM�Z��C[ďѱ��M��Lk/��������6�cjf���&&�g�ɒ�Xo9/2T�L&��56�_��W��̳�˅�R��^>WMRB)Z6��,���d�hbN=��.�kX{�ո�]+�j��3�GGċ{'p���@��V�F�<#���J�+�{���4i���ڒ6��E� 9�U�\�1?������.NN���,6�>fw�B4��5�Ȭ5����.2ش1��P���&u>�4=�0Sy�8�u:�4KU4
%4s��ݟ��G����؎_��౧������m��.�>ah`���~j�A7vl���?�i\� ^{���駰w|_x�a�2�?�'J��׿����;o��b�����h�Ӎ݆�HHT�L��?�\݊�XO<}�^��;HF�#��t�����薽#/r%������PM���؄�����������(���r��d������=������0����)�C{[H���U<��c�x��P
���߽{�8��I~�f��"�Fy��v�ѩS����7h�Z����ܜFY�J�H�=X^\ҟ|�i��Y�؆��#����ϡ���fkǹ�s�xm.?zv�7ڇ�L�rN��(�mDG�L���9MՍU$f�Q�������4ʅu�����N:y�:R0�@���� V�[�9S�*���jy�ڔ<�q�I�R`��q��q�s�F���R|C��b��Vr&y���G�j?��`>����2%Z_�yP�}(��ߋ�<�iڬ=�Rc`UE�9}3����|K�*.x�Q��Q#�d�#�K��X2%+�d<�P�]E.�k��#�ފ�'%��� ��(?���H7�V�P�r���$��`'���M�/�/h8���P�,c�A�
��������"�����..5,&�r,
�],�(Tr*VH'	�]��������7V"�~�ȖST�%Q�Xܚ ��k��e�3�!ڣal��s�r�^w�R�v�܊��ʏ�ut��p"`�0��x�k��B&a�<l�d�H[3�,nYl��Lyp��X����'w�º��i��r̨J����4�+���2A��fW3�恮1�=mҌ�#���&��e@�y0R��p��_�$�^Ŗ����;b)�9a*j��� IcT�G�:*��������}U���>:�.cqע�m!�,@DH��;'U�ㄏ=\�YdQ�BC�|D��1H!jň�I�W�u�b���L��G�6��!ѕ��"e�k(i�K�]3�i�v��&ʜ*I�c��a��M6�'��ze�*h�L/���<5�p`�)bn:������E��k䔏�:<n�����FE͏�eqM��L�d�T@�φ�)%:�Ҩ� �����P�Q�c����rW+����*��Zʩ�IX5CN�x��vƿs�m�'K�?Y�3�ȼFi>���M�5i�e=�D��|�k�� ![!;0O��o �"BL>o�RpmQ[W�3&�9-���V|��|t�8���ہﾃ>�}d67�a*2D�!h�p��sp�)L^��ܵY�������V�P�~�aY��
�0��6F'��5�ϫYf3�t``��^�8�1��䏰��p9bX^K�g8�n	Lh��XkѬ�4��0atw�~��;5eތ�h�N�	���(�����/:���v1����_~�s ܨVL#+�H�V�l�9yf�X�*T�B�n��xր��b	��٬��#=x�+�G�p?�]<��{NڜA����;�هB[8��W��g�W8}�*��"�U� �L�āM{�&�����>�(B�6����x���155�}?m�Y�S�S�Ŧ������%���OE�]*��z�&NSz�E�pG����n��b`[7�C�,گL���27 � \��|�l��.?4����0&$�
�r��ӀK4G�Rm`ys�O|�+�K�03�kKkȗ������4�嵧s^!��l�j����,V+�1�MUz�޴�u隩�^>Ӆ
�X��{�>��_������� ��_{w�{?|��g׎qt��p��G�o�^��ʋ���{FC^��㋟�4��F���8�����7�,��'ψ}`�u��^8wQ��ޞ.�`Y��8uS�A��ՎLŊ�xO��$�?�
�g��͢��1���<9sx�ؚ��瑘:�Bl(��RO�Z��Ƅb�<�~X\�C���r�p٫���αA�㺃�ePF�T`#��?�����{߾}�.���Q�0y�gϞ��Ғ6鲜Nr:8����هP$��9���BcFFw�KNf�����8�<*y�����:�l�( J:5����$�;�P��p��<Ws�em�y ��A,r,Zm��Λ
v�-Ah�T���������֮^�a��c(���(�`�V����I�N�
2eS@>#|���������ٝ~��!X�D.j�:�8x�m���kB���4�2��q��P�8�_q��%^&��mQQ�lE/b��aB6.�Z����@�\�B^�;-ȉ����e�����.�A0d2�R1���H�_�#����Z�����s��P@��)�M<�$���\G�W�q	a�&LC���\)���(�Vvr���Q�d���G�qw�4��2��rLlv;e1�@&�6�܊HE����t7	n~|�`����;
`Ea���׉h��ɏ`X["�A6[�0�V��T��dS E�B��2�]�-�)`�i�>4ԃ�C��<u�����²��t�ry|:89Q�iLd<���9���œ���Z2͇����%rdj	�~�"B��ovg
)��zո��2z�I&N�Bj��l��~��tR�i�(�g�JjK��x��d1O�}u{�f�r�L�8�Y�h�D�`Y#��7�����D~m�3��SP�,�=�'���|���r���}��$]�UQNjV��)Sj�F��@�&=�6�6�(�I�r��r	e$��|�E"�L/ͫ�&���8Q�V�kgS��+*��Y(�n�F�E��Ċ��'��n�G�l�PG�()��hI��բM��.I�cXe�4�ݪe�`���,��`qu����Ph�#oQ
8=�c�K�X3m
["A,�f��:pϒ�d�p�4P�Z-K�
sY�f	�BM:t�Ot��{p�|��j.�)�-^Sԓ�%��J:8�!��HnO�G�Zw�iq��&����7#6�N���h�� �쁎m6��Q��x�Q��g>���o�A&z�oi8wO��TP#a�#��y�KY9�:�����{�B|}����~|J����û�`��7����s���g�ѬҶ�
G�.�WgЇ�#B��y�%�ϑ>E��k��A��AM�y��Fw!�މ�'N����rP8��Q��-/��o�I#2��A��A���ۇ�t�*d���l�U�X�    IDAT,5�SIsY��qO/�n*����ݳg.L�?|��^QC�Y�;��6W�o��������E��tr$2�j�Yd3Y�bG6We
��G���������܋/�{�{�1�
ػ��x�_GOw7.����w��#S&0T�3�i4����sa���*��������܅�x��������@'-<��8Q��?�گ90�A��MN�\�v�ȦXg0�)���'?��v+U��1����h,"�H!�+ɱ*���⒞��f�U'p
PB1o���'댎�vtwv�>�-2�]���
ɡ<_a.K+�q|t�2^z�L.��Ɲ�3u_
��<��ې{"�	�E5�;^k�EF��}�M4I�e�U�j�\/T���*����'��_��_�������ɹ�O��;�wl>u�}���?��x��p����}{��/<"�������\�����pߐ
�t����qJ:?��`&��١|#.���݁<�N�+I੿��~����G�D!R�����EE�i~�MAze��KȬ]E#?T��5
,M���5���0Fv����\�Z��طs�=]ؽs\�"�T��Sb�������D7��k�҉[���]�ũ -@ҿdB0�1���9=�>,^*�I��^�F,�D*�l&���^l�1�H(,i �r���Kk���.b��t'O]��F�C{P,�p��<fW2��#��G�;f7��R��-´F�҃P��F��k����֮^�3����C���r�!OI��F��Jcg�D��k�<�������"���ARH=� ^;:;��ϗ���q��[q�C��tc��2ż���t 6�QW�[��G�A������I3�_����J�߬!�K�Ҩ�A��u{��ak&~|;�f���4�GV�b��,Z%�S�K�|~�#�}8r�������b��E�%S�EK��Έ���"�U�c�����/T����K�&��� o��Q�&G�>�[�0d��������/�Qk�����/d5! M��hY���Ul�'��gu�8���3�J"g<dt�K���s[����v(�F�6�D��ȥ8jO�w�`\�(R����j<H�"�k�
�	`t;��{�t]����A�)�dpi1�^mp�_����+�Ӌ\�����@���ϠɊ�'oW��ƝJ(m�y�$�E1$�Ă��IS�RAN<�2���̉(����O�2-~*�<�#ѩ�1�/�Q��[bv>�*VC�QB��E�YR o:q��gC��
� ���
�f��3C�D�nO@��5�ԏ�X��DץF����ynMH��u�ف�5lN�b�����'B�*d�K�E>;�p���� �+R�v ����W�;(�e��3�7��-� �,������?߈�M!J���V�9���C��]j���;YgM��}S�,�8�<`%k2	�
�.���S2��e���k~��
�z!'_�#���6�M&��״��ϡJ�"��e�؝��������Ӏ[�Ϫ�J��u��m,b�I�]ᤌ,�Rh�`�B4fY wcN@T�4��܈�4q/�d��1?S�S�2	�a��J��5t<��-���q3!�Ur���\���:��]���i5V	�h���7�+_�2�G�ceisS׌�����`P^韛�V�XMbuae
�9ղ4�'��iG4�Go7�Z�o��*56n�[q6FL�us�hw�ޏ��D8Ԏ��/����'��A���f3(Pצ�+r�yQ���³��d>{����nVq*����%#��4�NƑJ%Dg�n���B��nGov�:���cx��	���8w���ܚi�7�#Q�Y��X�S���y>�_�9I���;A	j[��������O�{������.�	LMNcdhXxc���o~�w��Եu��w�/��:��!�������r����'���o��o⡇��:yu
�?�~��O�����
H�B`� ���F�N��STA����,��vR1����dp��~�s�����(�~����9	�I���
X]����<�ԸٜbeLO^C.�F�M<����z��M�������3'���]���AWO�r-BA꼀ٕ>8}Sk�<����F����=�C�S�ZD��7�B�N_@��|��L����=i����tG���R�l�r��?��~��?�2!��k�|���bjv���X?�����n�.������go�_Ѕ���?|���/邞8u���p��>i�.M"y�b�.i~f�͘
ː?�p8d6-�Uvَl���������<�M��L9���%Z�o6^Z�XRIc}�
+�Ȯ^E37g��FAM��Lv�6!o��{btl�l4S�l��w���;��o�W\/>�D|��?�>�~�i9r���g���@�N4F�YP��v,/t� >�<��������6�ql�cr:��6��]����)T2�ʢ�)�k��:X�����ꡠ�lza�ki�<LA,���E�/g�
�cp�u�l��z6�a�	��L��kޤ��Ө�+Ed7W����%���E!��F~h�d���EQ=�q[$R xh�3��J2��A���B�@;F�Ɛ�䱞�a�����A3��Z*�D~��F�Ƶ�F�vډѓ�v�䐷�:���3�����eiV�� ����ۺ����!�R��,,�����A��J;.��K��3E��*����6��8�Ѻ����!䜼X��!ξ\T�e�P��_[���S�[\� nK��Q*�lDT�ܒ�R� 赡+�C{ă��z���\F��$eڠ��:��2Ւ��j�&���D"��K
H�k����ʱ�#z!z�(R�J��kBkX8��k"g��p5�ť�������t�(��FG�'9ldrB~��r��uF�ķe��煿���� �pHD�5:���nHd��)���"���O��1t�X.�������p3�5���?Z�Y����iW��"W�b!/jC������!C����˽"
a-�@&[��a�r������	6�>$_ȠXN����}�ެp$otQ�r���;Ȥ[����I����fF��1��^"]����_HgQ(WP����>u{���c��|��(�OL����{�L����7�SK4ɕ�+Y�=FwG��K^N�H�Z^[��i+����PD:������A~���ɥƇ���%�'b�f��i*[HG1�����.� :�P<�&K���<�j$)$�)��h{��f��͍c|�m`J����uN��K���@�m����#]��߱�bR-'	nPc�Y�����!�T6�������+�GZO�����u��l��� 0�e,�I�C��sM���j�WT^G8���w��+�Q��������%ңx�
�
t��Q�����}A7f�|����$cJyeQbͦ&7�~N�(R���^_�^���~|���d�i�4�;��L���.�����<��	BU�O�P�q�[�-FI�ΥSp;���B��C&|�*�6��"J� ?�5dN�R���\^ �e��rhp�g�H�Rǵ��h�$,�ޑ�$�ͥ[�1����?f�  �M�����at��#�Ƶ�9,���G=���"ړ�����${6�f�e�S(��|J�ti�hSD��H�L��p�O�������c7�ǵ�%<�����[��ge�Ix�.|��_���܇d&�������g^@�lR6y/y��Z���Ƿ��-џ	�||�,^y�U���I���!Q�j�E1��f>Ӗ�֩�����(��pYq�-7��i�ph�4� �-Q��q��5����X�'�c�Oj�������Sѥ��#HG��O�*0�!
?oq�@�T(�؎q�ݿ;�G1�}7=��H
�&2�r�������ƻ'O����*���)A$�:����"��.��!��� h: �%�a���<m5�\�r�M���7������4��[������x�}w�k��#_��.V�3x�W1�4-�W.��!\���0~��q��g�"ab|��
��4�n��vb���,gg�C�ɀ�Ć�M��/�t��?x��dӨ�o��0�	#Í}6��6�f5����HΞGi�*P\j	Xjy�)�O�������oCãh��l��Ã���q��>Y�Tk<�{�<�ԓB�����q�]w��r��L�yZ��`'֊���%x�.���s�qmzR8�|@��6D;��nS�J��M���s��?�LGL���F����f��N���2���t�D�wD�!{0�z��J!�P9�a�H���ZB9�Bfi��e��)s� ��̎n�93wD���;��&�ո��Ł��<���&yJ���m�3��I�!8��{Py�J�t��DZA�؈N

9�F���ل�m�.l�}�7��r���:��c�PƷ�IQ.V�2ʦ���M[�g�i�B"ml��>أP��p�U6��ӂ�`9m�|��� ���0��뛅7��d�f��"�T�%�`��� �a\��dS9�������ͥƆ�fY�Y��{hy5l��5��5T��Mߘ3�H��Gg09��J���M�dl
��ӕ��kC���'�O�^�PF�֜��t���̦7�#�l��I̮��H���TJD��L�Ѩ�f,��EoWD�!����D@[�߬�ǑLet��E�n��ZL6��B����+W�v�W§�����o��(I��l5��2Fj��,w�:R�M���ub�	l��Ŋ�I.�D�L�Ħ�T�XX�D*A]	���>ن�!|�
�.���>��x��w�4V}�r�jV���h�&-����?�=+_�N�k
@K�p ۶��V�������d���̆�� ����O��F-��L�j����סtꚖ��tqJ![D�J0�=���c�{��}�=���'�X���
��һ��bc0���k3��}w8iqj�Nx� ����Ζ�g��n�Y�ժ��c��ƛ�S#��<z�;�w�n=��Gs/����{����̼x�ܛ��z!�O�A����l�+���bp��a �/�����fF��&�MR�H�2Ϲv�G�4��X4�V�<�R9�Ξ(���������z�-M��`T�ܴ#���3��nNh�c`#�h��2O0t'�$�VV+�2�v��RCZ��9�{�,�9h�*r(<1�iB!_��Q�ytx�� 6so=�4���}�36&+q^�D2�D6�d6�*�*�>�)P[��rA`���6�|�Ql@��]o�3��8wu
3KKX؈�V���р�#������C�y�pl���t3A��I��Y �ꑠ�t͖iVԿp
K=�^���5�Ɛ���v���i�F��JǴ֕�S΋ۿE��}3��Zg�W�1t�2璦.������{õF�	;R�A~�ڢ�ɜ�֪py��E&��TI{�CN�YDk�4��|�_���o(/cfn�����*�ں	P�'���ǿ��7�������?E1�9�]��S'��Rf��z�ȗƃ~J�6A�w�y�s3s�H��2i�T�&�7 ��WL��s����ͦ6��Xp�7���,����FM\S��YXF�a���><s�t�\�1
	���2���C�熇��\�xj)81cC���VJ�y�r4'ڦ�ɍ��g\�<��<v��s����=�Z�:p��)���W��VKe03;�B�, ����֜.x��#�<�q6�e6V�����ojʨ�!�q�S�����/��П�����>��o��o���g��GF����t(�7�w��ӅJx�������*�m���B*я�����~�$q��BXN/�V�כx��8~bu{|�m�e�jl���Dpt?�y(�*!�6��+��9�@2�٪�!P����^Hm�������(�"!;��f|���X�,�f]H���s�=��>������4&&&4�f�QM���-v{%���mzn��˺�]]�'cXY_�Ȕ{:G�p�@P�%rω�p��7��#��Ҧ288���D����`��q��5|t�
�WR��ic�7ڏ`�v$�Q��X3#�V�޲�d�B�b�BRL�\�A��5X�)4�����b185�iN�H$u ���䴽D���FOW�l8��
��v�>p7�-Q19�B�[�{E}�p#e��5u�-����{j���}����>�Hw� ��Awԋ�C���+��Z�"�-a~)�W�ˣA��,K��;(Yt�Q���(>�E:�0������Jj�Q(�j��3�.�Y��� �F(�/��o}�S����J����w�)lK�+{�q�]�HfrL"�����@&WF"�G�^C��!dVtE����b�k��]ũ��X������
H�F�o$��`o�Ý��A�i���|�|	M�hAghl y躉�Y��X	g�\��ʚ���GA����VB$�Ǝ�^�w" �C>�ս�F;��z�L�d��g��^N�X8�����|i����?��܊��.�_#Yyfۍ��P�-�9�`��D��a�d���&
٤���Fp�!�F����H}r;��;���^~���N�ås��������`�a�M6m���ׂ�;�q`�x<f9_��D�d�p=�~��3/#�䨼��GE�Â��^��9��n6i���07��ɹ⩢\`(����-{Bf9��o��㶠��c��6�
�����S��]A*�Ք��%����mlC1GCj��'݌NlQ8h�KD� R��6S�]XD2�E�\����<�gx<a8��36ׄ��l�1��eP�
R��D/�]�14 zD(�W�5*��Y��C���FK+�XYO�Mf�����$�q��}�/� �)94.YF�Λ�OQ�5NY����e�beQ�������|6�tbU�]�!��vhm��#�@,�����
N��67Ә�O�nʙ�nC�#���0��U�;\��H[ u������6~ �f�����D|#�x��	�^9�\�9���1s�}\y�5L����n�ݪI6i~�L
�l�TR�����_�LOg3X[_Q���m��;OR-�b1,s�V.#U(�zA?�R�,�h�lX<���s�!���|�hXI���CrVZv�O29��a��d+hR|}6N���T���DZi2,�9�k�rp�=Ғ9)���a�l[��n�8Q+�Sc,�Z�@|M| 辣` ��
U�.�*�Ղ�2֔�J��Ki�<��ሦ\l��q�I0cea��/�{���g����Y�W�.�?z	��>��T�k8v�]������ݓ?��x�mĖ��ޒWȓ�UCg>q��
n�e�ۍ�W'��K/���?D2������ݑ�sch�N�䖳�F,<W�����1�}׭8�{����*�����S�29����l�B��4��y��64 '3�iD�>�N5��s�!$�"����y.HA*$R�	B+���@)�Mt����#�3�7��#;�F��O/�puj���6�y�$66�� ��{� :-�I��X�4�0�٢����i��
��j�ݲ���ˏ��W��.��x��o�l��?y����{ꩿ�H�n���{�����3Vݖh�F~t�ld�s]��������[!��r���d�YoW=�n��F�wwh�Ǯ�/�Y�����vc9��x�)m����0���ǩ��R�\�*���&O����j�D�[[6Ov�OBW�d92ف������S�ނ�n�Ai���XX��w��x���dz��w�U�A,�����'���O�D�@�˫��������qÍ������5iH��%��[�ƴe/W�0���l:/����\ n�D$�"���F�̔��'05��d��� ވ��Ӌ�<��@����nm��m�R@|v��/ �H �/��iЫ��Y:J(��x	K�k���Q�Tatkp�`��T��ay�W�6�?v3n|��v�o,k�D��.N �#��+q���VS#b���5VXj�V~J�L=x��    IDAT�F��w3��۷��ÚJ6W���&>:}����PR:soW}�m��Vz��S#"9tC*PH��G��!��HA>+�H$���(z�"���J��$l����ά��W��F��`t �_�.YvG�Rmnv����}��R�Kk%֨��!�	�(�v�B�RF$l��۱o|ȰKn$��Ss�:����8<
���:��`�H/�yL!�*ԑ*�P��R�F�d�B��0������z:����X�eష)h���:Ρ�+�B{���ٳ�cC�����@KM�ኳYX�X�4�a>X���X/L�8&��t{�0T�����@G�V �PFw����r��T.��D��C�سk� ��8�l�i#ɉ�>��sPx�����9��8�Ņ�%+\� �mm*��0d{�c����ؽc m>�4\+jd�m��M-�)��3i4�^:13����U	�����$�iS3��8"a��	�J���L�o O��ƟA�#8�#V��V5iE:�~�����3�@��`f:���U�?)��v�F�p��>�8�O7�O��Y>�jdN���&��<��`Qǐ%��XR�/��x
��r>/n5-�5�i|��7�(��Po��`h[��(�g�W�젡�7ܗ��*|�嚳/`~i�+XZ�T�G�
�E;1gi&%��K��kĐ�n9��Nѯ�����J�J[�g�PBwg;Ƿ+�gD���94j��HY�4��D"�SggpmjIϬ����.�&uH4o���27��CC��E��\���K��8��E��XX��ZC�ŒbG��+oæɵ�RG�^2����k�Us��G>���w���e
j�i7J�)!���:����c��5))���xO�|۬�n�O��Ӵ;QmZ�-�����x��/;K��R�f��d��kѸ�W|g��[�5����8<;H'�Q*"�J��d���4�V�h$�tg�,+y�9�M���ێbd��T�#���Im�r�K�E 5ԣ��-�q�tH�B�̜�w4&��A���@+��M\���ȰQH�Ӊ|�"[�k���j��><��~���w�8^}�E�,^S&Ӿ[n��o��]p�������3�1�����ؽ�����~��Oj��6�n���
�>�Ʒ������`׮	�it�y���x��gq��G�	r?���P�-j]��l�Z��%QV�"���=�Cw��3$�bz�2~��ϰ����D��6�f�`�-J��UÃ}��hG���c��4��}N�؄s�xܤ�D�,����2����5McSϠ2Z�WJ�*8Ь������#8v�n��&t�w���V��;�ěo��ǧ�#�Y@����.�'�Ȗh��S�)T&���V5�b�!(�P/2���Z.Q���CO|�k��{�0�={|��<��o���G��ݏ���	���i�w���(vn�X�ş~�?����������A3��51�ߋ�����92iT��Iڐj�t/�6�E��W����+�e�p��DQ"�A�#��EH]N�uؚ%�g������PZ�)X[��������w����E	{�g�0��p��
?�b9^][]�_��_��?�7܀щZhD/���ܴrH������\����uو�sy-�cw܆D"&A������ |� �$V�64rB^)#c0�+����w�����`6D�PE�f�z<���1��k���P����=E�T5q���C+>
��k��^~��z��i�^<�f.Ҳ��9i�æ�Qc�Ƒ)�kt�u�z$ʥ�o�"�as�e'��)�����>�����'�w�0�N{LS��C�T��tYxj}���Y��ㆀ"⭆���n���e���ƀf	�Q/���ػk}�a��t�������~��6s��11��j c����/4��b�@��`�d���{�w����r��ZelO�B7Z��6��������d3�u�㧯�ęS���Ѱ�P�1v���)�-E�tc�� �AjS�8ـ��}'N����3H$J�l��Q
��Ò�}�Cp٭Hnn�5��e||qsk99>P�M���G_��va�H���ЧLق\�<����Q.�v;�sZ4ዴG��Ӆx���/Lbzq��^O �ZI�ug�O���n�Y�yϗ���X�4��V��4E��-q���M��/#_$u�g��V�ֺ��*0�)�b�t����F���ń2	l��>W���ct�;Ǉ1� jri!�Sk�Â{�qY3�sU�ry+��ep��$�;}���xPj9u8�N����6�v!����M�:)N�F!�Z�l�jHgJp��X�e��M�.�I�ka ґC�p`�6Ж�B[���U\���ܥYĒ9��t}I��s��$���h�����.tw���vY�3Q) W'1=��X"gP�FE�{�{��T��kDd�f=�I��L+�$�I��l�t�"�a���&.L�c�\�<iv�Dձ���@*�S5:�2zB�݁p���955���Q�E1?��l����.��t)�$м��Ç�Ƶ�x�a��>�N՘� ¥�*�D���ЄL�`�N��I�att�aJ�I�&�[�
�����Of#��8�H�H�{�#��h ��_�l�t�6��g�+U7S���������P\\k_�(��,�
K@�Q�gi�ubQM���2p���^3TR��J�F��"�3�q��~�Kc����U�=��,R#t�z��m��p{�p��B*�x��6T���p���{�����pz<���aw��0��'���&gP-����!�4�{&{��譄u�ʤ�㚑��p�a���E[5+&O�{
��h�(~��X���h&��S�MD��O���c�qY��A����R*�%l�0-}5�$p�`���"�u7'�l�9(X[p�����IlX�M�F�&;��ٜX����o��/����ѱm ��ˏ��{�mX]^��?��_~��\���������ؽ�:||v��c��
%�r�P-ep�Λ��~�[23y�����s/ ��A.��#���w߁�>�����_6�;���+�aan	�no@���VNIrw4�rԡŨÊ�^����r="!��^>��^y	�\�Zl�`��rJ#hJ��]�j��v{m/���Ōhsl��v���E�7?�.sm"6��e5����q7ds\�xs�K��d���ie���cc��֣x��{18ԧ{W)Wq��4~���|~���{qqvk�J<�9K���aU(�?� :�!��^d3PD-�,���#���/~���7������Ϟ�����}����W�d���m���hқ�)m�[���k����N��#��Sx�ݏ�+��d���v&箧��{�>�3!G�r!��ϭDN����D�T����z��\/�v�+%xC]�s�g�K/�fM�Mh�W�:�QF[���&���;���fa�V�ޛrB��S����(�"Q!)��z�!�꣏`�D?Ƭ[c���E<���p��8�cccz�Ñ6���B�Q������4V�V����10Ǒ�ƑKtte�JՒ��N�%7��Ga����qj���,������Do���B()D����z�?�V�(�� W����텷�ug@(�l
��FQ)tV�4ds�>u�˗Dfkҝ'�&�yX�UY�jR`"bM���&��-JST���vо�#%Z��uȢ�g(�#�݅��%�+��Ϲ��r�lu�|���CdGX5v��B"ԫƇ�E��u$�k�{��� �a'F��`�?��ύ,Gtu�&���!6��% ���!.��h?z;B���So
�[�L*񒖥�T�Ix��Ƶ���0 o܁�?4��G� [���UP��x�ͬ����G*�"�Z/��ӈl8�k�����0K�O'g���{�13G����7�6&_���Lal{'n8�}��XY�ǵ'���¹�eX�~x�4d�����n�th'z�L�m��!Q��z�ҵY,��JL�ඔ16L�_��E\~:�Tq��%\���B�h�_��{�w�F{�&{���Z�l������xV����������>���G#���e��5#ԓ���P9�8Vx�L�cWWqfmT�9%Y�ڻ#C�URB�-MN��X_M����=��49�/�-��c~ur/��B�-�V�MC ��´U;�n�PW��t8ԫp#�*$���ėד)Q�(<�%��_X�f<m&d�M8,�56�lp��	rk�9+.M-�����k�+�v��v�4�����ng���D�M��\�.����"R�Q3dA�oí7�8�F/~�.;5PK�"[�m*�?�((en�[��RU��{������Z�R"�|Á�ë��o�.p��j!���;���M���AjKC	��#g^Aӊx,��)�? DЌ�-�>i�D�X�gV0��,7�T����t^BgM~XŴ>d5-�*�SOѩ&LAm5
*�*E�cJ�����{|HS=�������F�P*�~�m2O	!�c��c��KǦ S�����:>��<N���b͊�h��}5�-���6��s�ggcE��dO�ik+�ݼz!�
ڴ�L`�L��MpH'�c� W=�@��^��Oމ��X���O��>���q�l&H�����ɄY��VЙK�k�(g,�Bܿ)l�yO1/')�Ѯ^0��.f�s�Hl&Q�0ܐŴI�%��i1�?�u�
ɲY6�Ee�h<%�zS�|�W>34�P^J�r����q�������c�F.�B�V�Ή�x�K�áC{����JZ'�4Y�p��y\h��dS�ߣfQ�ԑ�pT_����&d����z�K<��r��{���d��B�"3������B����������~%K�kul�Vq�����+���E��8>:sO��\��E�aA&�Dqs	7�q3~�w�7�=n|�O��<����<v�V|�_�ѣGE�d�P�T�����^{/��
&�Έ>�F�v��c�0;�	 �s�����e0�s���_�m�݄pЇb1���Y����p���&�j�᠘������t�͸��!��e�4wH�TLkO�A���%s�(СKnc��h <l�N����%`-������$E,�%���B���,�_zq���������h����8��9����p��Q��և�����ƳJ@�E}x	�UE�$�,��r�X[�B7��}�u�����_�����=��O�|���Ñ8m^��<x@7��X�;�M�i-�p"M.a:��G�#�U�x��H�uv���qQ6\�|N�Z���ф�v�+6̮�pq����0�T��e܈�Vʚ�J��C�h�	C��4����O�t�}�Jq�k%��[����Z��Z-�!G����Q�-7��|�8�oHE����"N�8�^xN��c�;�s�N5lJ�l�8!�����
f&�Z��2򥢊�={v���:$g�g�P1����#��
[���g�N�������?�O~�Sr����Y,.��w�v�����S����P&��B��D��m}۱�-�n���P$mF�ldD��T�k��͹��a�d`A�z�z�&��+�!h�qn5�b�_n�ː]"W��[�<Z��_�;��\�ɻq����s4��NЖ7��Z"�H����\&��	�_��-��64	C�P�"�����D�ߊm�m�F[ȧ܇r݂��,�=y���XM�n���H/ڃN�}��M�nD�K�,����d��K"Y������e3�Z;wta��6���4w�C��[aq�p����݅
��v��i�]u�m�¡�D}N�H%�6��T�����ӓ�6�F�	�/
��#j�b9�����0&F1����/�,`�8��E\�Y�U��ZNc�7��vb�0���2�+%||�2.O��}�(@�50�ƞ����D�y SK����EL��>�n���A�C]*<{:��jdl��Μ�ćg.a#���δh��E����#j�g������q�D���p���C���D9��5)h�
*��6�,�l�v���C����&���@�l��b���+W�����w�Б=�t���{��P�Z099���\F*SVC@ABY8��M��5��b|��z���VI\�_��\�8n�*B3��fڅ�'�9��	��$K�f�K�پ�h9�(�[��K��q�!C�2\�\u,&�Z�#�\Cw���T�L�7Ӛ�n��m�|y��_���z	��vp�����@9�1s�Gڅ��9�l�kO�t�U���@ c�#r��R<�)W�C62y\]Xŕ�8���!��^�*XkE�R	x��!���~�\ �N+\���	*������D���!���� ��CƉ&�zqiW��b3����u5V�7Y��A����� 5:�ְ�R0�# u	p�N*uX&Fq�7 r#����ր�E6�.����^Ęp���nk�6����G��z�iO6���+�x��)L/���py�$F�tܰ�/��i����\���40R��Ǹ�!��V��I�H7_)�M
n%O-���ߍ��=���9��̏��s���y[��g�� ��`@\b>{DO��r��Y岀W�F!��|6�6�>:	z5����,Ъ%�R/�4H{#�LH�m�ݜQ���Ĝ��ݫ9(W��Ӟ�׍Șnk:GZ�:�Ɏ�Z�rV��{�������;;T/�I�i!�<��:���L5f�p�]U��lv��	�d-�{h2�g��n��{\N���و�bҮc�<���S�������.����U3ڒ�KgI��f&��=�US���x�ױ��!�B:�D-��[�����B����}�1��'/jB>�k����q��T,�q(�.�̹Kx��8w�.^��x�����H洄�i1,����i$�_!�A��|�ˏ����}�]X[_3�p��ill����T��@(���vD�AXmu,,N!����c��ppG��P͚�zIS}�at76��PE�&i���`�ت3ج9j�A=�6�*
t"�,c~j�.�`��`j���.|�/ad�:=��$��k����Y\�gqm9�,�-�S�G45�s�0Жu,oM�Z�dlJ�X��;?��_����3!�/?zu�w��w�b�����VڇRDC�x;�I +㚉q�ᨌ�]�gYo��q�Ѓ.#L>r`���j(�s�j���N�Z'b9���\�)��B	�k�*�����F��  ������7�yS��
k� pPhS/
�`V�6�f�'�?��w����MGvb��CӐK���_���,��:��?t��-/�"�LH��Chb�NY�}|�,��`sEj5��#
L���f���!�$wF��H$�<=5��s�-������L���{`e#���]X�����?��;H��>�|���9���<;��"�H �c�IJ�MY�(_(�\>��u:��UG˒,+�)@�H�"@d�.����;�;a'�鞞����^=�_����a�n� 
؝�y�����󼇛wV`ּ0L�P#��"�;��dVR���+�Q�\����f�H�z��F1���*�[0U�f��b�[I�ݼ	��Р,��N��J*� 0�g���)�C�A#s-em���pW'�{�#8��=Ƞ�d!����/��P~��B��i+�s�5��V��!�F�SIj~)!�T�&z$�Fw" ��,�!NT��Сv9����团��L�5������D�d��Z���xd��V���A�e�B�߯\�,d�*'F	�R�=~�:6����^���"1�L�޻���^~{�
��� e�Ξ��^x-M8e�gF�ܜ[��o�����狡EJM��hYA�Kc�	A��=	���s{n��w�-5e�CbѪ�J^��+��!q!ShaymG��{��ٜ������	!%!�jS�B,B��h���F3���L:�=uGF����(�'�lP��vk��< �+�ܬ(x�**��Ŏ�X�A�A�n۳'��R�Zܶ��Si�����B�i���!@}��Q��MhZ���3s�61���=)��DF'�?�@�@��"=�p��m,,m����DD�Gy93R�s�
��`\D���=\����ʺ���^�l����N    IDATr�&(������z��PE#a�'Q�L���0�݁���1�m]2I�{������,4gPҝ)�bC@��~j��Q���F�`e�8��I�����|?$�ݶ����qx�W6�!pb���&�޸����n7\>���J�<;Ƈ�1؝�$S_CA��M�MV̯�ཛ3X�Nð���`%���Q�O�m���9<|nva!|&�]�˻�ާ�����llmK(���)R���^����yn�6����L�i�6,��Z3Poh*����M��,�)���ix���bah%�N�hZ��G<�?z\|m�\�REV��l����=�|2�p7��"=�qdd G�d�æ��00ugo�{�LwH6��-����h�ddn�H�S�����MY�X#ߛ�d����3A�Ԏ[Z�xQ�3��`؅W^�.���K��Z�)?�a>S��p+G?9V�aQ��w���SM��gsBK�9'�2-%آ�� ��[2��q���k�����HCc2��I��ө6 �H�̗�;6��0�����BTR�ڐ�Y�FB���G3����BCj�����U,��
YP�˪�p���o�iV�r>���Ri�,���8���(�~�)��Z�f9�*w8�)d�I��SO=�s�=�|��?� $@ۿ���w�����/9=|��	�ܔA��Y�+�P�����_ċ����޺�b����]�%�Q�%������ob���צ����xw=}���{�E:��SSwp��$�_���V�ԾJ27�{_68�A���A�+�7�Etw&�_��}�i��vb{wo��.\|�k�F����{D=Q�汻��b)�by݃��8Ѱ�Q3j�W�܀��/j�%�''�WaGe0G�/�v.k>��X�Q�̍� I,n8,<$��������Y���cur�H_��/㉇Ǚ��d������y?z�*V��`�r�Q��f7/�[�`��hi�b�uc0�6��=�ؙo}�>��������Է��'��N��~X��ɫ2��%	�13ʞ9 �n	�	��j�`���e�-W�F� ~�,N?���F$ٍ�2��UL8�v$�-\���k��X�i!_!�ϩ�����MREi���$���Xs�^�,߼ �v`5W��D׬�
��B�nҐ�S��`�hX��C����FgGX��}����w|>/�XB�P*���ƺ`�fE0���S(U ��zG�%��2�7�N!_ؗ�_
-�	�ݽ�G���B�ݹ3+��#G�bhd�l	޽��~	�x?W��օ뢍͕Z�io�]pz�����v!Snʕv�Lf���&�Ey"����A�����+	V��T�P[�^*@��>dn�qM��J�e���i������ώ�ge�����Ob����7*�!8h��CMnh14��dX&M\���$)1�bԣ�D�I?i4ʈ���
"�#t ���7��v�%�-���������qt��<x�Ps�����b��.M� Wb�V�ȔH��9��$�E�_)����Ã���X7:Cj���k�9�]���;b-��c�8s�F:�p[��4j�<k��1���W.\��N-�.W@%�����ZC�d�zU&��p #���ܘ���֞�j�mb!�	'���ja�S�h;�)�����I>?ߡx�%���DV�"J��m$����D��BhH'7������NF�k� �9n��eܘ����$C���PN�iz?�e�R=0a������Vp�2�Q^"�P�>3B�jgS�����K�5��Ãy� �\f�����g�rC8��_@��hFGz���Ogj��]���Y�lg`�xa����r�G|85ԍ��L���]Kg05����%є���CqTt����V8�.���|�y~���dCcHC�pߙ����d��2�r����%L�,�ڴ�3�C�8�b!��8>>�#����� 
UG:]D�d`y-��y~ߺ�mBA�4�}Q�&B|�`3�"S���%+�M{������dkz.'�^7���u�#�����]��W09���7��큍�lR�i�?t�?$�u�D����[ť+���lN� ���)yR���N����S��<'8���G| Ys������b3
)0�8RҪ��Y��p��B��et��%	�
y�x�C��A�L��`��L�;����`'��&C��E�)��Hx\V���{9N5�|��M��8�[3�R\p �).�9BIbc"�^�Xפ8⹠�僠��:'DVǢ�awj2J�/��~i6�zj�7��8����-���O��^�ì�染|�V�S��!��-�S��u�[-�9S�;��<(��<��X���s����"���_v6̗>�!2f+�C,�U� م6�p����r`���f��SPޣ�2xa�5�jv6M-1A3h���@��2nT���N��� f�����䦆����u^+N~{�#�ض���� �pz=�կ}�����8����>����ׂ���������SO=����D8����v~ ��d�W��O߼(�Ê^�����=<����O���8{��5L-T��4�<Ei�$�$�����.,#�)!�-����nq��D% � �4CjD5�]_��/����"a���ο��W.!��/�[�}�
~��'pϽg15}��:l����1/Z6V��f�I�����,�$1����HX%)6K����J����y�ܵ|�mĆ��t�i�tւH8�#���!��1yu/��m�\�F<އ��c���?��O��ܜYǿ��ą�wP��K`!�M�[n()�f*HZ݄f�B�A&Y{�����ڗ>�����7�}ϟ���g��N�Od�2�EG�Q�hs����ҬR��i΢��j��YYG�ێ�|���I<��Gp��149��D� J^B�T�L��«o�bi�����#]��N3���7�"R���ݨf�Z�#�q�w�B�[�f�����6���*��$��Y��D�1��a1��c�>6���ݝ	�:{�Luө^y�!�>}ZP�4g�ӫV��C&Z:^z�ٌ0�x��ú�7y9��b���^�>!Jx�P+�K�f�O�`/���1x|�u���9�ý�H1=���d	K�{��J6?|�.t�l����h��m'o�,W���ds4���d�q���6Ѣ���4갘��B4�z]�9x���㝡.��:�BT���M�XX���N��g��ч�C�(c3�+��T9��@�~�!hO{���	X[S.�<r�e
�6R���tC�0���m���+�C,�Dg<(�}6*Â��.�S�Ǎ�ہ�ׂ�#�8{b>��9��ؔM�Zƅ�o��dl�����
X�����"3��8v�_���nT��(�`}{ْ.�Q��Q������pld�/���\4�p�������b7� !��w��+X�"n�R���>		P��|U�g�0Y�r�`��%��hHi�N�^�.�@N���K�K����9p[�����u���5l����̪|�fGHz����^i��"p���&t�6�x��ܼ���/�ԲБ�Fy�.�8��T��l���0��۫`��qH@��<;ju 
�6\J>������G_W{����֨Ѹ�>ɂ�:޿>�듋��2!��]��p��r33�hY�����iI���q:d�mE�Ǉ���BN&��Z��4n�-ana�|�>w-�U&�:�9�*|�I����l�O��S�3>܋X�+^)�xߚ���o"[n���@
�jA���9��D�Y�6�܄�]���N�JyJE�;F���"~'4)����jX��b~uW�2�*�~����u�iZ5$b89>,�W���_`s��w�M�Ɲ�Jy�a	ecրQ�!���N�V�O�.�!R���O`�X�?���R���!��*��:��ctd@��_|CW�7d+E*��6�(�����������[2�Pmv����1TzUbk�tG��G%�$_*A'��j��掐^�6����ϑ����1�˰(2�?r�)�<6�X�'w[�,,'qkzI�/*�&,4	�� M�j�*�6�1�0c��iؘp8�b�P�{��۴9)�ـ�:��Z��^��Ҁ��í�o#��H׸l}��a!H���;�F��1�$��g1�L�L��?���q��-?���D��0�7ᦀ93t�S�(�児�	�V��? �T5�K�6���%����6ى������46-2L��A��U�����Y?�k4U�6e(ԄĂ����ϱ%nh��`cv �:HNgax��Q�7��h�x�j�?�ǉ���ï�_����������o��E"%q#�C�GG,����82�޾Nh�d4[XZ^���i,�m ������r|�G�K��Y�t��YgX&� U���`ye�_������X�E>_�Q��.���r%�R��&\��^�����"��������5��%_��7_õ�kHg�������qA�ӬMi�������	V�j��@��D����$9���ﬨ	Hlk�����p%���Aؠ��<�4��!>P!�h���h�������5�J����*^|�U\9]�>�̳�§?����Ȕ�����y���/�f�C7ȷ�ׅR�.@604�Qd�[�����V��j6Y�����7����~�d�χ��_��������dw{��� ��Ύ�VFݠdH�҅�D+�Pl*}�*l5ͅz���� ������P_�t�,��B4�Z�unΧ��˓Xܨ�藆�+O���G�)"�<�x	֕O�i���6�ckaFy(���b��e<�g&P"B!���q��3,h=�����.z�;�=����J2��h��_ 	��^��E�ϩ*u١PL>RȺeC������r�ǉp������u���W�
Nq�i�$���`8�����lզ�+�XXNc7U<��ȁ�{��7��\Y�jE���&������^7��i9/�z1���J�h���F0�5^�A�
�;u�������*L�k��͠j��^4��!x���ч��n����Z�<*�z��!eZ�0����� x�v}���� eRn������v������ݬPYV6�3����C8<څJ{�j�"�'r��x{o\�o��`\
h��H8��$�er�,N�Za�
�EC���̤%� ](c��Rs��H�MՑ�>���1ĊX2�+]N\�u?~�

JJ�{9e*� �V����⡠�I%���"��24��ί�ki���d���\�����!��x�n;:�L��!���s"����t����-��,�gi��$��nm��O��,a|�[<DE����4WS�K�z��9X~x�4�I��t�����h�=s Z�v��X�Mc���?k$y65Ѭ�P����0�B�Z�լ�h�rn�Vq��&n�����fg�Q�F���A�@�!![�lW&�1=���ހ�OskN��#�����Ah��v�����0�����5�%ɥ�J��N,?��<8�e�KzIS�3�3'��bn ����F;%���?�f��q��-���p�Ip�K���x�':�θ6^k5���sxo�li~��S�y��ѡ>��t����hՉ�4���ǝ�u�,mI��DŤ*�_�eb'�U����=����F������XO�`���|���h8}�����iB6���ܸ��+��(75�Ba)�9��/>�R7���������J����l�o���.%���3%��&��LuE���e�!��""9��MhJC`55P/�e^ۉ�~���vI�Spm./�R\�:���s���h��d^��"�$M����Ȥ�;�x���q�p7�hg ���.~�d*���2�2a����ቲUYN��ٍEC�g%��9[8�IK�R�f	N��
�P�Y��o�(�d[�s9�A1�t3'����64��"mg(��j�Y��L�4>Ϛ�^��L��Sn��b���p�/���;`�@�Zp&�>����{f�ʟ��˵�|Gm�����|�"2Ez��ז&�BW����)�#e&�o�O�������H��5�7�����puϵ���I]t��{df(Xa6K_��W��/�/����?�3��V�@h�כU�E8T�c�>�s�ߋ@�/D��.S~s��Oa;E�_]�Ň��d��)0��m��2�ze/��-�g��AVf�,$/�vYx�ڣ��ܰ�sXѐASz� ����~gO
���{p��5$�)������`����D��"q#�B]+��(A��(�K�<=�bN�|��m�o��������;Ndk-Ec��{�`>3A3�φJ�*Y���\z=a�!x1h�b~j?|�'�~y!g ���g��O~�@'�����?{&����e����bC��Ca�`n�`���XB=�����_��|�D��G�?�������/��'�?�ć�K���Dj�h�!�
����uW|fI+e�"V�Q�T�@����c5��H�d&@[�-x(��&�[2��|/�6���:�.�,�n�qe��6���0��f1r].`s�:�'/�YJ�(�`�e�*%	�0x_X5��a�s��=]��E��+ԡ�8�O~�Y�vv��Bo���ޒ�bnL���"�!)��"�vv�L�J��p���yD6ņ���D<�!ʐ<^X8108�Pz|\��m�*i�g�37�L��@�S�AK�i\�\��V[I�j����� ���C�XE���fE8�b�\����I�!6&��"�B��u�6`��톀�/]$
��SIJ�r�|ß���uR�]�1�U��H��g��a'�%F��^<�ܓ;w�z{;���pXE���A���h���F��0RU�}���߄�"U9	ꎋlȦь�4����Ltg6��-�����='��3���E���ֽ��~��e�#px�"��"'�⁠Q��~C��><.�.�<#<±�<�wuB�H,�@Ѝ�ׄ��C�(b>�z�h�L���vy�޼+XY�9��C*�Js̓,ld�+R�X5!qp�}��gA"�]�)01�Y������~1?"�A/�A����vj�=��յ	�"��LluZ��܇V�bXn���a7[��A$&Q�7�� ��M���h�*�ߡ��!/DfV(U�$�� ��nH��b�q�+Zd�-l�,�?����b�#�
�������L}z}A��r�$�mu���ۘ[�E�cj�9ģ>�+�I��U�9 Zӫצ0y{�Z]&�I���gp�7�V>+=��Ŧ	�J.H&�@�W��. �) S(K�S����	M3�M�.���� ���f�k��X/���R5^��[���u۩�K�}ܐr���G9���S�^,������ǵ�u��4▆���٨��p�Ό�'�E�XDS7!�ӱ���;��X�L���u�,Zl&�2e��uvM�����0��{��fӐJWq��m1䕫fج^as�D�؃'���`u(�-�N�bק�p��*��� l�vP�M|$:n��f���:q���z�173��Y	��;�2�㦐D)�b�^�ʪ!��Ŭ	�efaؐ�ܪ)�Ǌ3GFq����L���	-�6i޿9���hN��Jnm�e�6h�5d����1>֏��A�;�(�,-n �oH��Do�����Υ b��$�$�4uZ�*�@�~pN��B���j�I�;'�,Λ(s0�
�4t�=X�����h��pY��ᆋA�-��K�7@����L�Y���4�ag�k����Kx��?�$Ų�:7c�M��O],W$�@V�1;��l��)bӬ��k|ǕY�@Fx0�� %��{B�J��m���-�L�	I��y�(���f��>U ��/T ��P�H�N��*�u�&`���E�	��ZJb�3� ��[�2f�f���>e�5�����K_��+���o}��d�bvXPmV�)������/����7~���Mt)�d[�TdyQ����}�v��2�����?~?�����+���R5�3��    IDAT��סY�0Z�I�S����'��k��4���1��g�ů���dj`��ܸ9���5��U�|nDQ�A�������@��C��|��=hXjh��(1���$�\V�����M�ڰ��)�x���->�J�G��1��������l ��0À��.������ayn?��˸v�*����������z�'/ /����'�3��I���D��vC@.=��>������_���|�X׺*d�~�����������9��O|���~�ӈ+p�$ �CUjJe{��]� �D\�'fs?�Fڹ9���[�(ds�y���q��'XUÊ�BW��A0�Mfcia��.q�7Y�rE�&j�!z8���8l�^�.l�\���;0W����s)r)�xP�l���(k2� ��tX����������c���w���V�p�u��6177'�Ξn�a)VcM�]��ueE����:]V�vv�;�"����OG� ��4P���dm'��YGW���l�YZč�Y즋�[�.���<3LX��K��4](ևS�L��A��$��zE6n7	!�sw٬��
(���Z]FugMi�qh���.e���(���̦�/�2x-h�����%�P�ŉL��<�1x�8��<�3i�Tr��U7�Kj���	�P5��o'�<��u���62�2n��a$"�:,��i4�ڭ������n��\7��;���.�Bn��N�1Q�Pj���x�'�`u�����?�*js�*4��^�rp#����h��.�.#�˵��:�5��:z�!�F���»_K���\��e0�"!NMa��sapͩ��I��|fɈ禌+Y1�x�RS6�^U	b�"*춋T�#�E<ꃋ�%�Zykܺ����cs;�+�/��������*#�40���P�Lj�5��^����i�;�<-x�״���R�U��֎�Y���8E��r�E'���.&)��s��􇐌�٤��Hn�O�P)��aaXڑ�N�%p���2�rzBXZ�Ǜ��ܗ 7��Z17N@Og>J_4�4�l޿6���T�u%;^����Ν�HĦt�Ōxjf�����v�6�@!�B�RG�Z��KJ��vӨ45�H{���*�t���X�%� �j�^�j�6S9L�Y��ZR���vNo��(`���=t����{��n'K��WEx�!%�J[g���h7�H�`X%���lV�9��<!8]�x�0,�Zv[K<(�c=�i@j
��l7n�a�β��l��86��S�݋��@�Z��E)[[�2��Zč�U�f1(�̔4G��;5�����v���0�>/V�WE�L��&yf�L0]��6~�l�H�t;��n�	Kd���w�3��q���85�@���9�mn���l�1���;K�QvdqJ�?D�̀@��6Q�g�T��#�0�ad2,�]�Ѳ ��㑆@B�^�2��Ɇ����[m��A,+Cq����&��9(	{Kd*����
�������6s���L���C�;ͅP4&hO������b�ڔ�����5��	;�fWk*��r"�����1����I�H�:n�W��~�܉LGɞ�p�B� G@L�jcȉ=,�?�W�>+d�k#BEn	��.Y8&�;���l��jC������C~�2x�(mj�YA.�TK�Y�pe�B"�Wάhp��M&���92LM�!���v6��F-�_����_��H��y�}|��~��t:?���A?���'ŵ��1�ׅo��_Cg�l;+���O�UT5��UQ&P�Q,a���$1����x��Rh��:�����
���fBI�D�%6�a��8rr��?����CG��p����q�*�FvB&e�4��$���KHv���;G(⇍�o�/�@��@�M?�lL N2 $��5
�H��猍@[r ���_��a���Z�(���攻��
�Ll:�l\5����.�\<���t��7~c#g�ÿy�������6��Ț�$3nø!�ĩ�l�AOX��Zn���s~�_���|����GC�O��7�������=1��ǟ�֬��������REBk8m$ݡ�-�II�jECg�[�J�R��K����#?,y9!�u^��s't^2yS��x��7�МQ1gP7kjT�Iި�f4�K礁�?1����ܾ#�������\J�uihdke\5��v;�:6܅�}�	;:��ߏJ�$]8��<�I�����y�֐��p��Л�]����)��e�n���Tj�lZ&����gN�������7�4�-�N���:*5R_�x��ܺ����$��5*��F�l�+%�A�AI��j���B\i�&,]g������{)l��#���Fr�Bh�5˩7Sa��69�~�"TSf�H#�S���Y7�ϏR�%?4 �u�s�������V!�L�(/g�ȕ$�H,jL2��j�D�e@�x�L�Ĵi6�ed4a�Z�AN�]�B��C|���=�H �]��U\�3���e��?;ћ��#��`g~��^����#��W��{7���O�
��Ϧ�U�ܸ�M��gC��%�,�@��{���`h�S��z�*��]R�u��p��R��v	�(�_��fo�w[y�\AXܤǰ0�a��o�JY����eij�����.A)�P+W�;����\�38�	��@��BW4��nI[����4��� I)��1�������Y���n�����C}���4���V�^��:�YJ�8q�����9f0IV��u�{y�v�ʤ)1Ι�qM^V��լɆ�t��Bv?�A���Ō%�d�a�Y����'�`�3��,h��uY]�,.,m����[�_ޕp=��?���(��A�u R�
Na��H����%]�����pb��!'�Zz�x<ChB��F:�wid�ƺ�i��:r�
�u���%�0���I��;e[��J����#���[9�������3�_ޔ�:I�m6$���?�8�Z�LCY��\��]��~�N�s�io)s�">��<z?�A��)�h̝�����l�����I2p5vj��	p����p��0F����ƱR60=���������pt0��>r�!�RV�M���}��2���l$\>�|�Y,�LVE�>�\A�T�m��M��� ��Saj(2�x��)=�.�g3ٻ͖'��6٩�ef[��If*�ڪ��5����C8�C�VF��-L�]����Hf��G:��A�L�Y�r�I=IR2٦Ο�|[��+�;��v�3�0���'��lr�˂�}���)�v~B�kû�N�h�U�!O��R�Ӭ�e5�h�SX�|���pR*ܤ�W�qcG�>�"90dQNz����Ҋ�w���>2�=��x���af	�`�[I�<�L4%7E�s�|6�_/	V��5~-2�����J6���+��k��
$K�N�g�Oj�P8_���ޮ� d�R�����������8a28�	rذ��%�nz��/��9��簋�:��*C��;d���%2?n�[��x����g�q��_�,���G�{���o��d�$���-��빧��>��݆��*�zG���s�y���"�p������F�(\zB4�T��3�D��^�O^~+�ۨ�L0D���%����H�݁Y��	pB��p��8��+_B�`B~�ć޽;+�a��5����Eܞ�B���/�Dw���p Vs58��ň����Lm\�`��l��.��| �����=�<#WlĈ�&��M�����hK��ŭ��O�e���#��i����0{{���0�N᧯^�K/_��t!]�:���l�d�҆f(@��n����{R/�T�y���|�+��w>�s�|����� �wh���SJ�ު��2��{p��i!P�r���������йζA����rZ$Q���x'���n�� ��� #���jMRtÁJӁ[s)����XX/@s�`u2����W]��q�*�حnx�N9��]�޾���@n��,��<X<`��E�Oi�������O���Cp;]��rr)pE��6�ړ������*\�1!S'^4^/Y��3r�[��l�H8(	�^�f��9���^�@9�p��,	�-TY�p�Ey,2�M�pub��u\�\��rJ�@��P �@G�THV�
2�,�������h�hH\�ɭm,�/ ��s.-�a���e<)B\���R@>Ѫs� ����ץ(�Nf?�%V<v��J��o�s����g@�^C�\�iN6_��@r&���͉2u��K��ߤ6�%���Y%X��?7l�4��&���.1fE�NxVa.;�v	���qg}sk���c1a�+��xHB��6���\0<�5`v1��߿��}I&< ��^r8mQh^{��p�������	ٌ|��\똼5#�mfb��ѡ.xm��0��&>>W�?x��+xj�h�l�[Z��h4JJ�f#��;�r��0����-%�c�5 I��9Q�l��&7�Q�ëݱN��J�kXT���&R5̨�[��X��ce#�t�
�n�����;SN���{���ݪ�}<p)��	�㦮Z��1�N�';V�w�<���/N`vi&+͖��I9�{nG�&ʺȑ��Rf�` �B�6H�rH!�qScn"�`t0���[��	�ש�5�by=�K����DV7�^?�VMd:D�����ʳĳ`s{�gW1��ښ���Ɔ�8��ȹ@2���^�2}.	y��H���*C�J͌��K�<1�L�,��:"-$��]Q/�z�"�
�MB"�aniM�X�˗ȗ����Q�=yB�++��M2,�8y{[�2�U�$уBS���<����XDg΂��37��1��)�Z3#����4�,~�$����&���H.��g�e.�cei�]��b�G $�'F�����$�XL�fn�o�K7��.ð��p�9�_����E�.u�ي�$Ц!
�y�/�|�Ď	�*j�hR����5b���`Qa����j�̼��܋A��K��Êýx��a٪2`�dwcaso�w�۰���yê!hQ��h3ͺ.K֊$��[�J-%�`��NL������ިF�@rr��+uO�Wá���*e5���Qk���-��J�<Wex�M�Zl߽�����c]ȥ�������HK8T�`QvK�x(�R��0�.��ϊ�R�X�9�n8�Ԫ,�lajzK˛����3�p3&]���ߓ�>���A��'�ɼ��P�V�	�����&��S�ln|�P��g U��Noo'��Hb)�-+��
Bѱil�O��3��Ѱ_h:3wnA�+�(�i�iW�L~�X)��C�9U��FP�(�7N��p��Ty>Rw����7~�x��GP�+x����O�}��z�y�|�ӟ�P"?��en[J��=��������S�ܥ_�d�Ѿn���J~���ە��ʦ�*���z����/���E��(�U:\���aS�ϧU㠉��z�x����y�˥���h��]�����zVB9Ý^��ek��(�$�<r�T$�_�Ī�i���,�=Rj��j��Ć��8L)kBVD
�������t.ލ�R����1Kj�>w>����v�/��>_��fU<�w�����@���IS���&{���x(�oq�M_[��f�'���o|����G��N�_��o�З���ċo^����v�iG�F�G���'?���n\x�<����He��%�GUΈA���8Wo-$�<��S�;��;�3848��'OH.��K2<��y��ݘ�I�7�qw�(&E��Z���z��V]&B|H$�Ns��`ѧ�\ˉ��MAy{�Z��t�l�x��?��`?N�:���.��:�~3�=pV�F�r�Y���ؽn����ЦT[�����c~~^�8��h)/�A:��ΞN|��:r~~�tZ��9�9u�`T�i�%��@�z3/*��Z)˺:����o�o�{�Տ��	8=��@�gu�_��&�3� u��h��x�F�B�hTudRIl��cc����lC��L��t��U���5m_:N���*��fv?�g>�9�C���hU�Ɇ�Ŝ:�����02���Vs�Q�N��U��4`mc��,�`c���������<ڭ��g�y8B�T��>�7�0���L�E��]��K�7ꃏ	�v���Yd� Y�*Ȅ���*�ޠ�l�Ĭ�-�M�\�<Hh u��l����فD",���s�e�W�&�q#�V�=�ΰ-��kEŽ�9�!x�wqmz�D?ܑ�$��Y/�U/�D�cL��ᥬV�r���=yl��J��(����B�`3��HL�:'3u��ή0z�b��IJ9��6����uT����GnU����v�3�kN�y8;�Π���q�\�AB��/�!�+lؙ2��^�ko]���&b��~U+"ܭ
��@8�B,��3�ٜH(��n?[���Y��b��A$�}G�	�ӄ�ǆH��ǁR���5�,cq#�������*�D�+�x�9-J�*��7qsj^�k]a���D���a����i�E1��_� ������4�C=��6&����*5�u�Zv\�<���I��VYE3��͐���k����;,R����/�
�2��I����Ӆ=� �!'*�*�
i*��y	�Z���v��˯���0�uil��$�^RW��!������]�Y�B�Bt�]?Y�)���<���]����0�����
K�/�X[���;7Q�p��z,83އN�ok�Y/�t�jXp���yi٪	�PL��rQp�񈡙��ĝ�������&�"rS�T(Ѥ���OE/���dg�AT]��8��u:0�ޓm����I��b 걡+h
WG� \!?�6���[q{~6�a�A��SV(�϶��  ��)9��ͳ�dsf�����*�x��Ta$�9�I�N�vC �kN��4͞I�,�ITAY�Hsۛ8���0���<�#ý�A[Y_���;�[\�~jO6�����R��*:>?���8�C#��E�z�
bP���e���-�2��o�/_|	�;��=�V���j�M�
#&���42����5.���8�� �:{�L����I�,�9��D�թ�αC�������H$��[^Z���VW6E
�-$?�H0�H8�B1���9	�c�֡���Y)�����ո�f�J*#�v&�����W�4��=��3�`:aK��H������{T|�צ��;/��_G���'�{
�|�i�9|>*���g�JY��i��޻���^�3����P�1<��C8v�d�L��	u���=]]���)�M����_��w��]��f�0ds��Qc=��� ����8S��Y��"���G��x%�/W����U�	:��$"'����4�+U���s�*���K< �?@L���@<��"��r��~�so��I�w	���^*�#�-Qa]�sE��,�+*�<?\6�����3���^@���݉卼dҰq�ei�(�2��B������F5�Va������o~勿�s�����ߟ��7.����v�;�07��jY�tE��g���z�����)��Wߕ��x� �-ME4��v�M���|����ƕ[��~'�������r%/锜s}N-|�i���4^zc�|q��>9�T��$W7��9��R�p��I FӨ�P�Y���$�'QJ.�lƺ3q�*R�@$�ϝ�Qj�qy�N�R�����/1�?���^�D���Yt��?/^D4�u/�gawθ�|�>���lll���,ҩ]���s���Ԅ�k�jM./o��,��8�E6�Y����-���7h��Q7�219|�� ��M�gh�2d�*�/�C��L�(�p:��Bg�J�)��R.�b2����M�`C�mU�c��C��	}�*_�����r�dC�9tAV�b#��qs�?��M�T�:��]�8�E�*�N��RGo5a�Dj���a	�Z	n�E�a���_�Ύ���{Bza�W*_�%    IDAT���Agȏ��wE�Z�JCL�4�ڱ�,���S�r�.\�(�ހ��(S�AC�(���y]v����N)V;bL_�粓����*�7�.�u)Rϝ:$�׊&xԑ@i�߹t7�6 G�jdZ���!��:�#N;+%5Mcs�ل��Ï�i�� ���
B�ir`!%vɶ熂27�n���Ɖ�#��G�7'��ݸs��!r6��L�'�дj�ԣ&l��0�S�2rE�f��Ҿh�]^���\�/�nbu#r�ܾ��_�l5j���튊.���|Ge�ca�d�L^�׻�+2}��x����슊|����s[��A	���4��Z��F-��$
�l���7���8�l�\��1;���yR9���=R�r+46�'[*���By��>V���/א���V��ǡ�^����R����'���n�^�N�ݰ˴Z��u v�������C���8���dSJҶv�E[��8F��$h�RR�J��ť5,��#�.���aw�d��kb�w������}29�3��)b��nͭ#_��`Ѹۜ�� 5)�(�1���&]1��bl��D����6�_�))��$�C�s��B�����R�]����Y4L^x"�T��Le�&"d%:�I1��ud�T 6@ɿ���FN:=dz�@��􆜑~�N6�� X�^m�yX�A�fT�ڑ{�4P/&��׍��!��Y���.c~ynoW@����B@a�5��LX�F�ŋ4<�9�m��=3dA&�b�A��LnUک��w�R�{�)�L�ą�K���"�cC�2��!8��g>��c�53��i�lobqe���"{"0����bA��7���phh��F{e��
n~��^Xq��\��߹�?y�y�n�Wʫd
M;� ��g�yp?Jդ��|�j��|N�1���!c``H����|��ߗ^n���ڐ�rp����O<�s�����͛�����vm�r�*jٰ����K�ڡC�8<>���~��.�����g�g�<��\��D���%��7�/���x�|�(fj������������Ҩ^�1���2�M�F$�7~����
�ɛX"Z�[9�2�X��ҕ��7���q��5ģQ=�U �x�i<��3�m�����		H|����G�BggB-�L�m�~�o}��v�$�D$���%���V�ۖ4u��ǃ���?���)yL��L�cm{v���0�a�7̎�BL7Mr#	��́`\�����`>n������h
IN�=��#F�9T�Q�7�js��za愜!l��Y'���f�m�`j0�ʅh ��H7n�|�G����%HRd�`�p�%�Y(��f�%e�¯��3��V9�Fa����|�W���sG~N6_�_�����7���LtۼQ9DMF�V^;>t�>���08؅�S�W��oq��|�"ݨ�*5.�����=�q����bki'ũcGEW���*�Op�&�U����񛷥!����a@�T���n�8iN�a�_X�aC�+�,��˲�L�݁�ߖ�B�E� �l ��z��̧$�~bjv���W����HD���"r�Q�O�P>�h<�9�z뭷�+�p��1�1)�Z�����b���$��,�t��#,���!�����Ԭ3JJŁA�����W/����2L� { �O�CG� s�r>�M���9���Ϥ� ��/�;���s�B	V�,����h30�ԊS��B�g�!u��喀���@3a��q|���Bl�i���tJ��5M�<`|�
Ѐ�0�L��.2���s!�tI0�L�`@pl�t�b^23�x0��-� �T�:Rْ��^�^�V:/SB�ӎ�xP��� �Z]hAV	@2��,��&qej�H�4��t5D+Z���ZY�W~�݉8�:B�����2�����˫k��	�T�-���NFWN= �wM���Z�ݘ�z� g0�7 [6����4��7[�d� S+�W�y8re�I ���Tq���I
"&��Ѧ9��d[�n���&yj���ǩ#C����4Y�X����w��ʉ��H~��!�Fw�)�����5�WӸy{	{���6�z��BmڄN�
ŪhWC������#���H�#vH�mC���Ε�%��d3��U��.ac')����^�&���l��ڀ��eʹ�����X��V��G��Ƃ6�G� ��drH����*�n�I(U�ER�!��D<�p�%�"��
{XX[�l�n��
��{0���'�q*==G��v�*�T���aG���a7�������iwV��ۘ�����4�qy_x��x�w����L�cquS(C�`�b4��*e�|1�vF�8qd�	7jzS�|����W1qkْ�'(����S�/���6�l3:��I�p@���ĭ\�:+�)nr(�:{x��B�G�'~&�x��MḼ����}Jo�@'�=B�%~l D�HiY�S�>l(3���Rn�֥���j���g�yh6C��1����P�_X�̣��tI�ު�{1>�-~S3�`�'��|�!�'�,0���%\{ɱI�R �ۍw��ҲcC��� y�%�r%�-	��ɭh[�d��!	Aj �麨V�m7<���
Z<O�ux@�����tx�x�0���Z��T6���M�R)ih��vwS��:lv���0Cx�6��A�[4�tVJ��˧aW�L����"R�y��r��m��-i��!
b=^�4"���=��U�"M��(c�����>n߾-�gJ���pX��!�o(�=r��s��˫�X\\��Դ4��NJؚ�)��Pȇ��.><����������<��{�m .:@ {'ER�DK�E�r/��L���dw���nf����8���;��[�eYV�,Q"%�^  :n��}���}A���svN���s$�p�}���-��y��vX`7١��pSL0;?_�i�dL��+�������7�~W��7`�V��G�����Ï�'[��O��ӿ�-ܡf�{�}ػgBV��[-��p��udstv�J�/���ׇ��� o=&�N��
}���}�Q|��F�X��?�#�:u�l�<���򻧧.�n`zj����׏be%&o6�,r9��-��e��m��i��F���C}���M,bauE5�p[ �v?�6=�.J�|�,�;��H��k`m3 )�BZ�wUC�s�-[!O3����,�~=�O|�g�9Ai�ZC �~kT1�J��6�����t&�5UE���49��n]��į~�:~��W�J�3�dC���b��h�|6M�m����HlZkjم�=���?~�?��4��߾��S�����1y�Q�s}>K-aܷ�s�<�^{�M|�;���|�H&jک5`p����������~����s6���&�5���7��8S1��d/�}�s�Ai/%p{-M���J�S��\�$/�_�bh����ZDtf��	d�3h�@9	�$X���áC���|	]==�11����0�yi����b��=]�p�.��U!WL,�9y���y155%]lww'��x1[PU����Q;�.n����s�㴡�+�Gy����.�<)� �po&�ǵ�Q�����׏!��
Ҫ��Q)�hݸw���3�_��l�����-�kfJ�D6�p?^�����(��H-."9>���^T3�H�@��φ��G϶�8��� ۨ#Ỷ�I��S�)�����M�C�N������*Bojo�5腓i�Z�z��cX^\A���^l�t�;F{[H�<��"������i��q��L[wn����V�,��a�Z@d�b<�������a���_Kcq���R�bV������<��-2�"W;�Jcbj�3�P�^椫���f�������,��z�z�M�^;v篍Cos�����Jæ�|�xJ8������DkGX
N��n-����ނ�x�D�
�M�l��g����Ј$��j�&�"�[�w� |N�0����-�8s�&�^�M!C�����{��ju��g��㖧a:�����b�eR1�l4���<,�۬y�k�x�'y���p�oB/���I��RL�2�����[��5pct
�#O��tώ�c��m�f�L�������x��(�r0X�r���I�w����k�b�`0��U,��|�&Ƨ��0Za��Q.S�O��v`��GTj�\NL�,H،�8��=-�}pڬ���M�j<%Ġ��e�*Iu����[��Z^��͛z���$�8,Hkaj��s�$���H�Ӂd*�D*#Zv�ށD:�م%��m�B����z>�~���CR����|P�֐���y����n=\���J�2�JE&a��g��o �6c�`�4-f��Ê\��I�<7*�)��#��-�طm@<�l�Y��p��(�O,��s��)Nۍ&!gq+���]��pBh��t�;��>��f���b���`$�,�k��:�Ӏ��?�`q�
Ҍ�x,�|.#�dܹe=6u�Í���Z�pȧc�Z�R,�R�([1�t99����2%yl
��,��Fn��D�c�(�F���j��%�-Z;�)������X�M�5}�I�,�F�r	c^��F��N�_���=X�ւ--FT
bɄȧ
�<���P�Z"���d!�Mxlu��/	�s;rngRi,/3���fRɜH�n����4������d��sa��p��G� �BIDJ���g-�4���/�r��lK4��ccks$���N�v�i"�4��H�����3>�FGg�=������R�8qM�2@�G�@t�r3T�E΢���wpuxL|K��/�����4�a��}�� ^~��q��q�݇��}Z�^�J���:�.N�:�T6�C��'>�	X���p?���8��i>0ȕ�_��gg��≧~���/"K�\*�������>�Q�ݻO6�\Z\�:��|����ѷś�&q�gJ2)��u�����&7�fG�]��k����
0"�O"_�Cg�#�ꅯ�������EE�ae���ѐ���PD8�ܮ���
G�v����m�O������_�"�%Y�!���D0�Z��p���sF�aҌ�f��*�J�K�����E�Ջ�ז�Ϳ�1�9>���a�:œ��q؀����GC@�BSqv�������?����c*����#?{���=���u�Uy�M��Ղu|��b��~��<����^��J�P�ٝ��u����ۺ��_���	<p�0vm�3�d��ë\Y*&�kfܜ��wƤ!�ٚd
���v��'��5<GU�5|�Q߀�mA=�Dry���K�d�P˭BWM�VL�a�?0��|�#صg�|���E�R��&/��;�������h,,yp�!��#/�B!'�,���H�adl�O���p�ho	!����K��;�J�;(*h�I� \��/���^9�d�"aXd[�$s�Ύ��~ ����JW�'h���,��\���4 ��x\q��q�����ͣp��!P8��͠��E�ʉ���ZC�A�j0zT3�j�V'�fv땊�4x���چ;z ��J����Cƴ�=�E�()����5�c8��ʍY�~Z���=܄����fIN�ԋ���."��\	�ဠd�[C�,�т�Dg/�alv��Uѣ�I��|C_���,�8M��S2�p����x��SH��"��p{|� p�N�k:�c�Ⱥ�[eZ�I���@�R���<Fǧ�L��4_)��q0��n����֩$[`�;E �ڱa;qQh;n_`--��Q�Zuz���F���b�*+��]���b��B��=l�Y�v�����8��-Y�mN�,�JaWGW؋ݛ�	����CF\����W�P��Z{%'�
�:��	 �w���h�"�R��ѳ8��E���~)[+-$��!PS���qMC�1ӄ��I��l��A�`�&-)Spq$ި�.�S��sW0��"[��c�z��� f6�`ԕE;y+�S��DΆ���tf��m��k�&��QR{O����(`bN�[�s�����B�lTQ,�t�s�iԨ�%�dC�a�:d��8բ��K�'q��$*��fu��D�Q.ee�?��C��=Z�������0|^�55�0���l� ��T19����8T�j�BAҐ�U�-:��$f���F~��H����*�]�"�M4�W�fT�\S+(�3p��R���Aw[lf�ה�4pad�{�ȇ�M~��l�iž���p�f�|1�d'�]å�3�г`q�$^�Ɯ�����DL�4����R�+��o���"|t�{��FD�-�C{�ґ�ԗ+��9]n!M�j&���.�q��5AS2����m�qh�D��^4���d��K��<2��X���n1�k����y�3K��g6颁�ba�����q&r��H_�{q-�MJ5	!7���vC �Q�$`�_X����Y���jT�4)p�k�M]Ctj-N#��*�v�Ж
��4���@���L�I�a���Kp��9�s�� �ER�fff�P��4���JB�?Y�(p�E_��)��Y�!�����!�)!U�0�k�QRDZT���x&�>�2h��2A8%#Ԃ!_V�:�[6d�"Zd0r�����ٍ��	\��B9�P؏�&�8��jÎM[���'�"��ԋqu�$.���XVp��8���'0<6-�,R�L./�n�)e��|�cl�0��W�����w�×��%����,��;'q��)���L>�<� ��/�f�/��:~��pmxTR�+�4j_����/}Aҋ���8��),��I>T�V�?Є��G��c��@�<��Kx��/���R�H5����g?�q�޻�ro}W�_@�% Ԡb%/hӺZ��[sT�=D0��0)�zL2P�ץ�A�mk�}�!�<$�g�h���
�Oz���`�zQ���[�%c��.H��'h�[�� y�Nk��6`C m)�F�B�0	i��?�3\V7�:C롯7���zO>�<�f4�^�6 tˠ�y�Tl&��G�IÎ
eh�|䑃O~哏�ׇ����&��_}���_<�]��Qm.�4Peq��J.����A|�Gv걺��o~�^��J(�A�0���G���!����qkr�uw�C:��h}5 �Ɋ�yj
�Y�����E.5�1+d�J�/u�l�	������H��=�9��ƠdW`��_G�)�-5�������؍��Rٸ�y�twvb��mp9�+jF�N��%��� �̈�v�4�*z��������Sr��ChmcrlW/^���}�܍�N�h�u��
ΜƯ�y�.�`%��7�O����h�k����0�ܘD<Q�8����/)=��U#֪q�4�x�R'��NQ�X�buz
j,!��$���,�i�&I�]�ZC �f>��i��7�D�Id�I�
�����{�!0�(4(2 ��;�r�/r�\hI�$�[�Va�D�@Dhg$�f�K~֚�.r�sK�|�V����;�zDjR�2���?we�t&/���,�t�=���qKک����!�C���W���A8ҁ��.�47�,��,�TY2�Ը�"��4�F�L���ctlF�����*�V=�A6�wJ�H�47D�����]Ǜ�OI��?�"�vJ��^�5�u�����P�W�p��A`��|^A��ex8������hAs��ф��e��Ob|��h�C֞�d�uu�����z�N
y"dPl�0����%)�t�:�z[�0�ĺ� 4�JCjE:���%}�jz;\L��4 �4�Ya��`!%�D�O&��JI|=\�:mF��6�����D�ߡ5A:�� jUZP(*�[����2V�I�9�=N��c}o����*���u������	�.fDUoԐˮ �d��wlA_���g#G~<Q��xWe*    IDAT�1��C5R�g�{��JN��a/tL"�qWH/��U.�����عm=�������[Ņk��y�@Q�6�mF�i�U���)��x0m۽FIF2������!��0	#{jv�G��Ӣ7{��9P&����zE6TNka�Mr�m@k��tK+)�Z����i���03��G�d.���*�^-���B{3ַEZ�vpU�G��������NH�:'�0����Chi��f�ߌL��c�.�&*UPaq��Pe�� !�N��Uy]��qᔸ"���6�߸�DT<_,"٨����َu��h�8�����A��BCW��!sV�l�Nn-6���S2�6!|���}[���C5��D�T���WnJC��q�i���b�I�+,>����"d�k��Kb��k���E~�,d9��3FH6U-���?�D�5,�y~ަ��t�C �7����7ZCE�����Z�F٥q��'0��X�y&ݯ�� �"��
�DA_ �]�v�}�F����{�5���sB���l�P_��w�bQ��Ή��Ɓ�ΈD.���Uԩ�2X��$���96/,f�bCj����|��->;j�,��P�yfp[Dꐃዒՠ�9��I�L��,��3�u�y\�aj��� �L!�� �N������8���	{�m�̎�l3�㵣V/��=�;v����	��f@B��3'�l���42�"&f����g/��T7����d������p�TH¢/�s�>�ǎ�'��g�*~�ۗj�����\��#�8��q���jlI��x�A|����v7~��/��s�����H�wQ��?����"ҙ~�̳xᥗQ̕Qa<�Zm���o�<��cطo�3���8v��z�)\�~]���C�җ����ӈ��i\��+�����%�I
ҕ o��]��Z��m����cA���|���|n3����6w��$ UkXgh?M��4���"a�}R�x������L�:7Ԣs�4��f�Ѐޠ��;u�L-F6��Q5!艠-4��o�x_�ۧ��Z�����mpka�N�	Tl�Mk�BI$�qv��|�˟����`�������g/����b�r��Z�/�ػk#���p��5�NNb�ƍ��G���N1t��c�t�:����+7G�/a`h ����ap#����`��}��g�v�N[L��UF�HZ�#�Zpu|o���|�
�3�1i4635���"��������� �"��3dE)�Qͬ �(�Js��4}:Tdr��F�� �{�^�{�]���2� a�r!��9U�f���!�!��\��x"!�/�f��a5;$`��9�/�N��]�����AM�¢d��y �}�.�v�DL�ȉ��O����\3�������"U�!�փ����c�֊�kD���/�#�����b4����\��O��n��y��e �jEi�����^�f����<b��$C�ܖ)�y״�lD�G�h1/��C�q��5�$#�՚�����!N4��h)��\M�I�#'g���:t�i�i��~���4�����Wp��9	�9x�4�L\)��'�-`|fc31����z�se���lj7���a��n!�XL��K,x�]��KWoHb���Co��!�:�bx��Ve���U��&F�����E*[����b��*J۷`��-"u��,�a���\�"�Q������U.�H!"]!�Oc�P�mְ݀]R�W���@u��p��u)�ns�y&��V�Hwu��f�Z ���gf1<>��ŘH`8���rh�qp���v�`�!��a|~��I�F��pꭖ�n®�}��l��a���hr�	���x��5dJX�~�1Q��TX3@j3M)�!�R��$2,�lx���pXL��]p��p8��;��@a4�Ɇb�&!X��X��9⮗��ƞ����T��崊�ct:�g�ca� ��J���upϡ����S�g@,���r�n�`5�ȶ�����=vA�R��τR5��UjZ��1LJ.��Adm�7���)[���U�<���(���80��:�~5�%�5�>��>(�o���E�V���� ��&��AscI�r&_��+7$8+���I��ʷ�%y�6`S�m�Eo�咦�^YI���IA�V������6���̔Y��MǱ��w�؂���I��ɩ�cs�x��i\�X���l3�&�4�X�;7���X-:�N��|GO��|4W��S&oܼ�P���BslNB���[׉��v��dB�*�ͫ�#hf��^��l��Gw((Ġb1��Mj�M09<Hd�ȗ��'��62)�ybt��~;܁��I��T1 S�E���lL��-nz���>]��A�T�\ �e)`Y��%	����L�e&�� �����4]�1A�� 0�hc�[iX�8��ɴTy��<�vH'�R�bת��U��%��8�+�(��V+hr��� ���P�U��U.+�)j0Ԍ�W�#;6�����w�!�][7bۆ��{��Ƥ�#���J*��3Ө[�*:,��"��ٹ�ヽ!�*RrZB<O����Bgw���&F.c��)Xem�@ο�+)1Ƭ�P��q���?@� �"�ŎhYA�4�jYd��o�c1�7܌��կ�����N�=��q��qXFX�FDZ[p`�l܈�p,F���VG�vZ�K�!(ab~���O�։p�[�o�'��Ãl:���q�%��
����h4jx��w��K�,6lَޞ.��/b��M�,. �\�R�`߁�x��'�7Z�~�_?��旅t����~᳟Ɨ��EdK��?��G�B1W��&�k"��?�ٵ����{�l����ַ����>�u��ԧ>�{����,��$�Vnaai�rV���R�lV�V�5nc-@;��AR��4�T/pj��'�qY�Q˯�h� ƭ���
�+<vE� �5����	�F���V�p~��� ;B(�k�P/9��֞��F�3ə+��/�^_D��aC�^DgJ��7�׎^E]���n:JY��}54dpɟӠ�I8�Zɠ�Z(?�ȝO|����i����=?��K�.���;ڠ3Q�a�G>����^x�E��������'?�!�`/Z���ҨR\���b�<p�A��<��[J�޻���A�|:�6ԉ�\;��	M��=��^C��7ɴ�:\-�Pk�v��r�@,�rX8r:̂�4	ư��Pz`V
(�o��^D��(�'�������V��䰣���'����< n'�<y�������s���%��7F���o���������dZK�t9PQ�_Y�j4*ɪ��I�7-�+��6˴cqi�8��GO���<�Ul�f��r}�7a��]0:}2垚[AMg����x�2������z���D=��Y���t�Eo� �����WQ_^�W4�Q�7�ZK-��V^+eN����pǃ�kA��|��vX2@�����^C`P(��x�Z����b}_����f�*����8m&d�u������;W��5B
�ɹ���
��H���������`]7C�X�8��������|i9�D*'>���>t47��)�^'I��	���)�K+1�����*�5�LmN���"1:v�vo���"ԤG2Z@*_�U����C:����-X�e�4!����1c��,и���bu��a�23՚�����m^���mp� c�S����)�y��E�Z��4��`w�{?���b)VXM�02=��sX�qC�09�z�-^��>�u�A�Ͱl�������x��e)�ހ&"��v��b�B�i>�xa�/�f,&+��<�p8A��%Xmӄr1+�xCt&!pXm��r�O�xk�;��앇�;�Ã��,�=}���"�@�R1�u�~�s����ü�T����E\�:��x	f�z�*?��P6�����1/F�ə\�2�|�*�D�ɈJ6.�����:)��Aob���R4�Sg��}n�d�N�u�b�f(�����m"_	5��T*ȧ��&㰚M�[����^c�K"s��
����*�!�5�Px�p��4Ў=�7 �Z���8C�N_��|f[ v�_��F�u]�J�ز�6n�ց>D�v�wч�̅������Dav4���Z,*������;�wkg;�cL�>q�"�o��h��hq��=W�m�#�ZA1EK��{�> �n'��: ����gp��E���8CD�֡!l������*t�����(���\�[����y)�MF��"�~�s���`uaJ��ͭ��8u���b8Y��Ch��Pt&1�k��<�k��K�d3�hkFGG�Hʦf�1��(?#	a�ru��5l<D&����FdN����L��X�	�H|Z%2���L)�j��i,��]Eq�t�$,,Y+#[*#Wִ�e	��&�,$��ߍ�®��11|��铰�뎽h���%�&O�nu����|"��K������f��!`Cύ<e��|����;=}w�q@R�o^>��ѳ�-��9�YBU�m%�פ��P�A�]�2���A�T+� R�%n#�ʊ��#�������׾���N�`\���7�b~iZ��`�	�6n���m���C0�f	��JPaz�J�B�|����_��Is��&yR�N�[�����g?�>���1���N�;?�1b94�u���Oe�YI �����I|���η��т_<�~��066!�S�z�M:|����t
?��S8v�42)n��y<P+���{������n����w�7XZY�y?��.8�F��sP@	p�RK�E��W�H'�/���s�cEMGJd	����0�V=2�l�6d=p�3��/@	1�^�2����NiYK�L(h
H�U��D��h�1���B �$�&��+���F����vj6�1#��m�{԰���@�v�y���o�?��Q��F�-n(�f��R\��󆀞�j��b�C���W>s��`��������ٳ߿5��>��ٍ��G��o}�{x�wG��7a]O'؉��v�]b�
�]�B4jF4�Ə�4�9<���~`PX�&���PL�:��5�x���l`i�a-�Q�Uu�CR���$�I�bQ{�B�VT>�Jv�~7)4U�D�ƲL>fǯa��48E�(]:-�ڵ��>���$^|�E����b���C����;q�}���r���w���c���hk�ȃ����N~��5�D&!���6��^U��eF~:�%��F����M�FT��W4�xL1ٰ�ni
��{s�
U6��S
;���YX3��͔ɪ��f��>��L)�P�I}��*&�_��J}u�m���������5�5�4�1��C"4U��`���)�P�\�W���#�ݚɕ�T�e*�'ΰ ���k� %=m���h�8����DF�	|4���|%��"t���(&oŐf�Q�꤀tX�����+yD�.��@OW���4C����f�X^��������!�^>N��ʠ&J{FL�.bv�dRLNXln(��T��`p���mEW�I&K�XU�i�M�g/������J\�P���mX^]�j�����ZqTfHW]��79��>�4[f�*䟽���uc ���r:)h��LV+�'�q��,�&� �44���؉�f�a�+We�2<qK���:i
F�x����D[�~]�lt�Q�)��ur���|� �!MB��q
�BF[k�D6���R�eBKEW$ѵ�w֨I�*`��d�\���u�&N��}]a�t�ć���Q�\�>���/ciyU���K�4Љ��6��9 ��b��J���Gp��)6.��X�
��ހ={���-�T��	�~�,n-Ť�qح(���j�����l��9T� Y$����qsbN<DLj�ё��)�tj-�.l۰m��}��[/�`ZK��a��X�I3p��5)���&�%��bF-3D�Q��m��C��l��e�89=��g�bx���^�/*�JI4�j�&��}۶��퀩Q��b�pĺ����$�<yc��pxCp9=(�pJ�����]��a��^@i1bnq	箌��M��8`��&ic��𺥡�R��g>ý�����/�Z^cD�}�4%�v�����҂��6��0�k��`&S���FFnAU9Qf�Kdz����l®��2��p��9,��Wf���3�_M��jt�{͆@t�hC�V3q��nۺ���XX.��눧3b�%���z}�\�7�L�g���[�n�I�X����U :i���<�}Fm�I�^��U�Of'`(&�_�A%����_SAe�R^K/�P��P�eii���z�A�ޱs��x�g?F!þ�[1��'^'N���l��ï3=���xK�,R�:bI,F�"1������u���j�"��-�v n���J���j���) [=_��t�X��T咖��T`3}'D^+
J'�5�RY��+�c����������8x�a�s\�.T��x�	c���Է	�P|,z��q�3LA.G<��P�B�82����BEo��D���r4)�j�����9���gç>�0��{�wx�����/��(
�<X�4*TJIɤ������׿.r�g�{�z�\^-���b��~���g���
�����ɳ�V5�����<���A1C����0>�ǰw�.��N��g�����G>�A���b~qzSu�;TmT�Χ1���X2&$���6؝v��E��::�[�)(�2��j���\ߒ�I?$��!n��<n-V��>�u�\�uŢ?��%��������e�p�()�uɦbc-�m��-׃�~ �׌�y�4�ZF���ܰ�c���e3:}���~���Ë�,fkB]1�nk��9��D�?��v6�J���<�o>��PC�w����|anu����{6��C�`��ܚYē?��h�9�t{����۷`]{��:e��v�5�?XU�I���1<x�Cضu�pQ��`�K>+5d��ks�!X�ՠ��a�:u7%Al�uB��g��d���2�J�Rf]^���R@l~��W��.��]� )GE�T�]�cϞ=B�x��$��\t⩜.��hq{���u�N�!1Hi���$y]��@�E��N�8�1B�J,�/cnn���+&'���bs�l���E��#��%ŀ��n�"�Pu4ff��$��h����5w�L��{h)���ee�V(1��m�IB����Go��{��=Բ�!�2�ְ��/ɐ���M��G�����.�)mp�n�{�~8#���!�M�5 5���I
0�>6�M���"��bY�֐ݭa�\vX�u	�bAϭob�ix}q@z%>�(dnW&gWK�`i��ϔp1�O�e�6��ٌ����8�6���xH���� ����|M�� ؈�3�Pd��^*��j"��xV�D�$q�Թ�l�`<���͂��0ښC��&ʔ�}��h�e�L�P)���у`ЇD*��6�� )�8="�J$�x��Y̯�`q�œCJ��QX��]X�.�� c�\O�:4����9:� &R2���5$�}��r�IܜZ���tV���s[H�#����6��+ ���Na�p���Q���E�F�A�Y*�e$hi������RR���
�D�y��/ѳ� ���-�j4���B:�g�l5x�z�v��܊`�.Iz�|n,G�8u�<.^�������9�����d�(���N]����8Q����ۣ���[�s{��ADS�_��q��0N_��L6'�M.�n���v�א5����?���(����RQD�H]�A�K�]zl�Fo�E�T4�qJ���9���<�=���	Asz0�d�V4��%Swkt���sK?z;�0�j(W��Z���ØY��h��$[_��2�>'z{:�*�
�N��Z^WA50�����c|.��P���,��ɨp6�w����r��F�����1�F�y���f�S��l�>�Ⱥ:Z����})YE&+�&�p��,�R�0��0�$lV4�U�i�SS��N&]�R7�j��V��	���bN��a'�o�BogMO�    IDAT^���;3�ɳ�F�.�`sd����1���I��E4�Y�fw�ڍ;��,���g%��Ave��IksJ��	���Lf1s�*�����Ќהn��]�Ezy��֝A���ʆ�ii�m�CI/ˆ@�ĥ!��V�tȗK"������
Ƶ9ģx���عu��c���?�č�������P��ܪh��0lr~�	dj
��ӋQ��.�LS��JU2b�	������!R�R����h������x��`�J�<U�ehztI�e(b�($*��
�7�\��مE\�>��7obfyV���o���=�L����I��|
��G��F�=��{�b��6!�x�>��6�I��t[U���$�T��k����������P.�٠��X,�dH-e���/��s�����Ͽ�_��e��>TUn�̣�cM���R�j�|��}���7����o^�/��-n����:]��bƟ��?ŧ�����Q�Rr����jE���U��R������%�r%���v`���h�'���/��ʧP��Q���$e0�{����(P�>Z�P�U$R1ijl�׈[��Y���b\�[E��L���!n'S�}2l%Q�>�/ZBa|>4�(�M��.M��O(���YN�iݠ�&�l��ƾ�fH���I���1���ч6�l��iބN��x� 0@Ͽ�����b�~8/*Uf��$��V6�A����ɮPL/��<����|����!������^;��R��im���߉?z� ���<I%7nB�7�j��Jӎ	�`]m\�:� ��TK�k ����ś��^@�ߌ����u� �jU��t�� [�����P���,�i��d���u�!�;�S5���s)Y�3��^��j-z�L�l�P�%��8���"�2��60z�HD��Er�A�/�Jo��,Hx�6������Q&�5񿩩Z(/:Ѭ��!��)�Q<�6�ml�;�����DĘ>#�:�� ӻ�j�#�!I���D:DD5�<,]M��<�Vƒ��N����5�$�Tu�0p�c� �Lcuq˳3Pb�����=ɐȿ�yQ4�(���ZL�x�^��0,!?��"
|����	W�Eqa���u_%c�r$�Æ�`���$=�M�niɅ�I�A60�(�ilt�*5A%.ǳ�ƙ[A4�󟞅���D*0rMHҒZ��iA$��;� <|X ��F�rr�@d�r��A�3��R�WO&QS���r�0l+[�����k�l@0�/M�N�	�z�%Ԍ�}��xQ�J�d
�L��P3����/_-������N_�]��o�uK�,~��H�1�\̠Z�	6���3kk( 2lJ��x��,�y��ӆ�21�����k��ZH
z�� ��+���f��X�H���"Lz��]*5������y�$ƍ�C�O��N*�ľ�Y��M��S���#DݴA�5 r��|��8	.�BB���{HJ��i�,�>���U��H�	f(dK�%������[���GxƵj5��\�*pk9!Z�T���'dM�#���C۱cKj����`P+n-�p��y�--�������a]W�'QU�V��[���k��R���l.��E��Ȇ؀��m �����ކ&za8��iF;�a�bY����8{i�*?#l6�ݥ�)9��ө�����&�$��js��\�1%�3����y�tvE�u�F��#�J#����M
�?�b�0<�h�o�U"�^A5�Ǒ�݅pЍL*
�ہ\���XR��<�LF|MAēix��D�m�zir�٤\#6��r���1<6��ފ*osru(q� ��mSI&�f�ր�I冉�%����[	���+�<��:,ܾ���׌;lG��%N��������\z�K08Q��~!��3�����bۮ=b�>w�*���ّ���Ĕ_��rI�-�)�v��v���L����L�g�4
ZF����<W�i��]��e�+�rl��`���Rl���[j��%i*���W���G?��~�#X�ہDto��"�&G1�ӎ};v�mwh0R|֊s�&r9�zT���f���-XZZB<��;�����Q/d���Bkg��
f�'P+���ej��i��,>9n�%qV�Zh7.y�t�a�a��P�V%�����q��y�����k��v<�ÌD&�w�ǋ��K���������@���*�)u�^HG�f$	1ٛ�.��~�s����g0���j!�Ɖ��A)WB��F{Њ����>��$Y}�~���`%]F:_B)S亁^�%�ri!�������o���^����J��%X�ZC���>��D���Sx��S�-����l�Zn�j(Y/�6U��F�ۿG}����,`�V �d~K47�rh�A��_��-GC� �:[`u�-�a��V�e��I����C7!Hմk�9<����Fx]n�<�B���d^_M.�N�ȅ�����-�����JA� 2J�(i���5�����3�:�o��KJ��d�S,p���ڀ��8sz
��o~��9nH]�����2����\������)�T<r��'��˟������	��_ki���211a�_�|���\�+�����������E��:�0)��ڧgՊ<����,<�v#�mb|���sϭ �)J�#����QJt�#F;
������Y�؜�5ê����W��!�Z �/���"2L����RD����C)��B�h�ULܸ����~��F��
�v�)M"�_�� ��&T�L��ɦ�]/C�Jfh89a�ՁwmK����f��)�,<��D����U�X��8'/�2`s�� Y�PK�F�$gs�#���QB�Dg �_#���g��bQ*o͸,���Z~�WT��]�!1?���P/��/�h7��bN�9!�x|�sڱ��>�8|t^V�y�(Z�Ь2��S(��9�G,�J�	Wn4☌2��V V���Do���.�	�r���Ax�L'ҹ��a�$
�\��|T��Ē� ޔN�@6�U�ߨ��PUbwb����2�߄;����˚(�5��FCb��%�r��{�S�t�(M��bL�Œ":h��O��bѕe�l�@������D�"2�d2!��j��	=.�
) 
��"I	3���8VSYxB��9���,j�4�J��o�6lܲ~�z��I1��بq���6 N���f���㝓�MW`uQl5�?C����[7u�����rb�BY'\��7����㚱�4�
=E�Z�߻��FLT�tr��;Ԕj1�Zc���?�QWE��V���L�Ђ�T��7�u�*yX�5�6c���t����\B�^-<b���!/>��&�l5c5U�)���Fg���aF �'��$3o�Ѝ�C=���(f�rM�+
�FfW��e%���5,�7&���N��.�,6�5����^��$Bs%N�4�>�m�䷷��a��\m�c�Faܗ�����3W02qWL6��e�	2_/�WnpQ�JQ�����M5I]��5���fB*����"��q����E�3��|]F����쉷�Fbvi	7'g1��F"���h�n�eb�*�"\��ܻC��s(Vs��aѦ�Hk��y��3E��_k����$9�����p{�҄S
6���� �)��O��P�$�D�I�yC�ٮQM`Ҷ7"a�GP���8��p����l�I~W�4���=3����y�/ŰMJ�¿�v�%�v��.��TJ�
��0�{|��%"=}(2[�������4;m�d�5b�ךh�9�`�πSv��T��VihR	���
�sN%�&wC-�jb�Z�*�	�2iJE)�\�	�%��0&��c��G���=�t�.�}�t;6mD{W�l|Q�s�f�g�P�4P��*7͕��(2��q��2��|���(�cHD���BC��Q�'`pjC5�s �5ɉ���&���=�Ao�����yx��//���x�7�֩S�_��lݳv��F'Ν�ӿ�)斦io��m[�~6�5A���	ה'����1��09��:�����\��bt�������w�����?�>���(��x���/~��Ÿ��T��ެrKdD��D�Vl���ݍ@�	ӷ�$D���ⳌF������'����|�&�s/��e���X�h�\�(�m?��@>�Dk[�~��8|x�x(r��N��,��0�0+y:��Z8��fu� �u�IN�R0*P�*��5�$N6�Ź����/)bZuI���M������s�.��nc7k�ɬ���i��ÊJwI���^K�1���R��[�p�G;�!�����W���h����y._Z��~���dP�[G�O�wX�C��635�ej9�jf���G=�������93��_�|�?��6�eWS��)���|���.��N�u�u�C�s1���|�zK�*�����UBH��X]����4�͓�;���0�6nl>��_���(�v�^��'A"ٵA��P �<��R�����e3��<״�\�il�*v��<���0#[���U��E!]kxJ���hw��-:��pK�$`N��C�U�.��0��L��e�bܲ�Hf1Ia�Ɓ�����X)��r=� ]*A1���B��FX�!��4�5P,�u0��|�đ�� ِ�@�iDr!+b>��n�Ĉc����$�,����4��*���ↀ�71d�/��g�φ�Jɐń��ޅ=��i�b&�^C $��V���b!(��rzY����Y'r�֨�<������j�C=��w�Jpv�8�"��X��ϔ�A(zon|$���̆I�Z�m@I#�k�UT�s��u;	�7����b�B��,v�3��Z�t���vx�MBhᦢTQ�!��Y@2�	�V^L6OW�,Mt$��=(��qM�׮i`�VN+��ɔ!�6d�y�W�XM�̂��D�TC�\��K?
ѳ�_�aP�b�f7�i�f��ȯ�P�����N�[��Đ�OI���L�(����s�(v�m>(Fʣ�0�*�$��,����ÏP�)��U��a�RҖr�2�6����E˼#b��υ�x$����IC�Y�A�\�]^H?��tF�����4W("�a��}�!�9]r�i%z�&�z�)Ud��m�ӋE\�9���UD�UPI��}L�IMp��)2�a˺v���1��V���CMBӌ(I�jȔ�[/�ՁZ̀��e\�8�h��M���ԙ�K]8e2�����w���;vnD�$3�.J-U�(��z�_�1��O]����b���y&[s"����M�ZEKЍM�:���e�	��Ny��$��%�%4�Y�Y�~���f�H�v�{|�U+��gg163�h����U�F�	�LE-f`�)0�d}W�q]�n��eF6�o%>&	�
@O$-�������@ZH�D\66ަ����L�5_�V�l�x�ː�c�͙�+�u]�Ǆ���\U�Ar��g8�����|���9BFڴ~\V�H�L̝ ��`�b4���[��mIx-�l�GO'|^R�*�p�0='6X�>�pQjDj��x����$��g�������ֆS�]��������`H97Bl�J��L�l�2J�u��(�����(�,6��L�T��0>�����AoG��".�9�z6�ݛ7���]�F*'���|V�9��G�PC����̒��׌6$�E��)�<voۀ�����쪮E���ԩ;�A $$� ��c�ql���66����k����d2"#I		P��[�թr�:9�{ǘkW|����]���Vuu�9{��֜c�p��T�do:��L�7R��  YZK��s��:mrCR��	#]x_�F����W�P��q��Q|���߹�C�����Ძ�]�ܨ��G��}�,�.bp�[��(a��[020�T$)��R���	���L4�Ӌ%|��w�އ�֡aA�j��N�ky�@o��W��/��R���W��o��K9�;�k�e'�gֹ�vMZ4�htw��.��߇��U�K��V�Z�/��f�|�-b#0����A1ϳ�붮5�)!'�y�!�3�+y\|�y��׼����%k�Ad�8>��O�@�����|�`(�3��Zڷo�2�={w��R�!�,PC����|�h�k&#�4d���@\��sH��Q;	���i�` $Bܐ%k"N@�l5z�2���7�&�V@�C���Ջ�R(��U2�f;�p�����;r!�?1�~�N>��Mt�M�7��@83��!�3����6/�w�'��G/������_?!���]�~�����Gސؒ�"$����p�۱{� :��Ɗ��G�&�	4C���A2-_��]����J+�yZ�����S~�/�EPjt�&1�P�7��}r
ɞ��$m������~�Pov���刔�cفM��(���?�Qi�PЋ��E�S�@O=�8ٽ8���p��C��~S���LB�� �(~�|0."��Av�1-�@4�y�6c�	7���\|������rŒ�C��ڦD�@��Cr�c;v!38�XW/���
�z�>G�I�|.�Z��B������Ի���*�T�&PxJ�f܋3s��� �"��&oB`\�_�X���KطC��a�.~=�+^Rp�����3_xZ�����PD�)
p��(�@�/{_@c<b�ۓX��5D��þ�"d���16ҏ/:W���0��E��3_�0���Z�nD�wEQ�������Э%� �`)k�JǑJ�{�A�\A�X��ڊ�;�;w�ęg�EWO��C6LDeNOLcjfAM�m~�RB�B���""VXy��7����ү����,�2�^,,�`e��we4k>��O�B'B�vn
z��kiR�j��4�{I��א�Ǳg����+ǂN<�T�uK�əe��A���Bj����c�0���4�ڹ�[��k]�+UL�,�#��T����E��,#�a�#��R*U���1�C�T��/��@)���D�n�� �0kN*���fӏj���"eӞG�^P�pO<�g_v9�{���RXJQ>kR��#�Vs�c���CǰRn(��k��'�PX\�Р�����Ͻ�
��1�[������P�D�H�v�@Z��ࡇ������
�z��P�h>��uk�;5��5�K/>]]�9�i�K�y��u���_���;4�H��F��Me��sE��Q��h[Fp�Y;d����T_�5�$�����%,��o�v$�|��l�j5DB$#)q��V��8��i�+���_�!�U�p��SA����0�ҡ\͕�:�̈́CZ��>�حTY�
�W�@��o�|��P����#���c*�c�^�q��4���=�9��x�Iu��}����s�#��Ѻ��"��G"TÖ�.��<$��K�twi��5�c%�Q��Z>��:`���'w����C��+��� U�Z�>M�Ho��uDg1;l¸g�[feK~<�9�����BH�yDku�=˚�H�`ڬ�Y�}r�]Ai�:�UĚe4
9��(�ٔ+�D|�r��
j۲m���|\��8c׈�~����,��½{q����Vf0}zB��&�g�&g�Pj�����q��Ќ�����0�}p�1\r�^\t�ػm��RFR�.Q*[�U4�g������3�v�h_�Ã�d�4����!����R3>9�o��'���~��-;��{\��g�P� _.�!�Ɲ_A����X?��8��@?{�0�?�L<�&�������/�F ��sE|�_���=�N�[9 ̋a�º���T��	�+_�䖗�}_�򝘚]V�&���I�b)T�uQ��8��u��tR��k�V�!�I;�w�^�ܹ[F�'籸X��bAZ:4�p�N�>j���c~a
O{����7�{�؂���X�. � �m�����iT�M�Lt�sV(�4�Ʈ�����-��uPiW�,���,=R���F�D؇0�L�f��ŹC�e"20�$iOʏյ5MX�|p�%l���lX�(L��"
p*��It%NФ?h*E���$x�=;    IDAT3�:5}�m8c�%x��)|�cw��x�e�hE����KVWc��ۄ�݄ ?_��W<�S�����s���X����~+���G�����n���ߘK%�{����W4�>&F(��(��hIK	������������ف[^�<�{~q�/�����Ϻ�[��{?y����|�Zl�s_�NLUˌ�IX��dKH��8�<��8�M#ZCݪ��*XTJ`j��5ڶM���V)���X$��t�v���ǱCG����y��˔/S�k�1܋�5zM�P�F3D�h������0�m��1Ca4��+1W�z�b�lX��G�=<��;���G����_�-���Ew����4��lz���r�j�,�Q��ksGB�N�	M:G�T���;uX^�	������Dym�]��#:�O<Z�����'P(�m.�'��|ޛ��b���y6�}�-���EI�^��^&�1��)W�FSv����D�D���(�������P��<����B%X�s�P��Hui]S�G����7����U,D�8Z�JKs�aAkF
��l��[���^��E��7���k)���_b����M1�+�h��S��曜h�tO��bll�#C���R�>M�����F .���CKU����)_�	^(��,�x������a�B��n��-�H&�[>77���YM\����
63���#h���,���<Ъ�ZE�<�yJ��29N����&u2�H\�;�� =����k��`����Xo�m��5��e,��\$�޹>[�?{PIǺ�������r+�4HD����e����޴@���ݦo��jk��C/�@4��?Lڮ����^ɪ@ٳ}W\r���%"Sh�Ȥ�Zi��bl���p��Je�ϸ4.��^���,��Ry�誔�N ��;���~��!���!�23Wŝ��f旐���i3\�����&`A?�&y�J����at���*рhr�!��I��5��I���g�S�B�M���)<��I	@��(ڝ r�
�nd�4�j�����zi�����k��3w����`d$f،��fgW�i�Po!ݝԳ��k(C"�����I84�t�H4� ��~��X�9��Ŵp�=Q�ׯ}�ɵw�ʖycM�B����I1�*�|t�;��b�����E�0g��dJK\���}��KE���q�}HT�'Q���	��
��h��'�v6�4-��g��T��:�''\+z��y��r�����D 5'Qq#���⌄�܏4����!���0/*���nz��x��W#��QX�S���O�/���lIw����J.���0`z���v�tE;vG&'Q#���Ș����d#�]8o�V�F����mx�}�q?�&Q+��E��P��|����ए{��9�ǰ`FcPߐH��\��%|���G�x�.���3�?�J	��xt����]_���i�{�Yؾ��#���8��$Z�G�F
F���7��?�Ǟ�­�~r�~b��,l�)�6�KS�>�����<�9W������{���;����U*t�4ې}R#E���HS���t
�v�/hw*���)܍�s���hu���W��k����J�!N�S���i<��k�xF�����a,���i��)bfi�(C�"	s��ҠK�R���k۶1�¼�YMF�4I��3ò�H�V���[�xJFV��c2q"�fneiYuid�D��>�,v~��E�0s�se��:�?��Ʊ:�V��݈`2!%֝�~2͛�>JR��X�}��8s��x��Sx߿'OP���K9�$��R����_�Sɦ���k��W��E���W��^}v��o�l��ߺ!���̻�?x��C��/��#8��~�L̠;��8��,!ߪ��fD�NA���l5+���n�
��W��[��_��6�+.��#;Qo0��iߐg�F��C#���d���>L�5�ي@4m�nr���ۑ@�OT����ʃ��,u87[Y��jS�j�R��A�� &���o�0:FW(e�8r� �<���(4�U�FQ|7n DU��|�8�Q.zң���+VE{a��!E��0gdr�;@���!l=��lA ����
�W�*��Lҟ���ܺe���Wy&��V���g�!�5�k`�į��8���	��-D�����)̟:���,|�\�\u~7K*�]�����j�f��ˣ�G�Qv�D�̵�<M.H^��(��q����Y/|��S��(�\H�����vGw��R��L��ZMt+�Ѷ�vݎ���Ƚ�겙 ���������MFu�
��	?x}i�G��l��_�͠�
xE(@$B�9�$�;��<�nb�#�(�C#�~�a��Ƈ�M��!*�ü���9΂���������'�Tʇ�l�؏ɩY�3�Ʋ!3��o}��b���Z��J���,{5>W~Dšg���KMEV.�S�`���#�8�3JNKI�~J5��$"A��t���p���ȗ+B�#Q�s*���^�{kٳo��z��oBn�zIk�~�΢T�+�s��Y
�/d�G�ߓ��F}��z�euH���+zݬ�ff0;��r<���V�

>l�]�i��B�{4J��v��
��Q H�b�Q'����c�g���&��lie�E�tsb8�z��Sۉ>1M�<�$���F14Ч"�rww7��'~�q�i�b����	�[]7ڮF¦C��)ãx��!�am�aRM�kei�R	
񍖢�,z|���p�z�\�s�X\^��V(��Xh�k���B*�h�L��P?
���%z�Uc�������4]]=�Jw�ȣ��t8"��(p��
���abzQ���$��қ��� ��xM������6��g��5h��Zm�f��c#����Y�v�����RQ�O:+��\�4`���P*��G������R�%ŏ�;�?W󦡙�Ϛ�4����:s6�ux���+�I_��_�]v���޹����h�_~ťi,O�DquA�2�P@��+X0�"�F��7�`2f?�Zu�?��?���q�jUlK��5�F-�&2M�� V;>�ZXi�pbf�,OJ��tm�]�v]�r��q��b�N�@���yg�Ǝ�ў�����V�ҍ��>��/�������N̓IT�ŒXk�q|y��?����ĹO&���wa��]�����������/k�u���c��]�P����;���QW��Ъ����Gw �=�pt�sY��c_�w~� *����C	�VZ���Ǟm��m������Kw�_�&��
:C(�%r���M��e҈��₾IﬖVѕ��}��%/�'��w��>��[XY��i	m�n�)�r�kK�I{�v����<��k�淾[��bbn�jZ����;���)��@�+�`��y�����M�R��NQ��q���_�d�P��ɰw�s���5�@"F�v�� z�z�5�=tmqqݎ��#����	Hq�6z&��s-�eC@#�H(3���6Z	II�F��H �X0	3�d�Q��\��<�~�K89YD�у�?�N����݅*����r��l�y��_�ꗿ��������[5����}���u߁Coݱ��ƛ��+݋;>N<y�==��"h���*83�P ���jL���K�v�=�R��w_������]�-��ܳ/���Ս�X'��V��$����ů��+>5�D�.�
-�NZV�I�Q�������B2�Kk�RUa:��'�A$�X�Z߷V�h�50<Ѝ�L7��Nڏ���xh 
0k9��(|$7���l���7���)��nK�3(8.� 7�t�]=�����g"��'�A���J��2�1�	�É����{���R�u�z��F��դ�!��+t
l��$���Cvy	s'N"w�4���Q,�����M��E�¦�h��G�+RGQ���@�=��`�a�m�\z�5������&��a���6<Є����tX���+�y]]� 	�|�M��tB�:���X!��
G�|}� �F�R���g�]�r�,ʴ�؄IX�`9���0$��M��ZԄ����j�/�YD�y�xp�@�3V��I�D�גMU�]r2�I�#�?S5~�(f�14<f(!�$�U�5�]�&N��cG���y%NxH��R��U���p2��>lj��Tij�|�Yҟ���
+"��s���W.&V�(�^k( _��A���gh�v#^�G^'�v�mt!7p�Ŝ�|*�%�tk���x>ּ�j��T���o��m���<��6�H��֝Cq�����D��AD�)M�x��Y�r���V�̄�h�(4SR����J&tٴ�n��Q��~�����~2��b�IoBE����d����N�V*�eu+*�\�8)�h���A��Ҋ�P�:P;@��E��+�Q�$����6�G��g�V4[L�>����L:�]�v`xhH��ם�ܫJ�V��8��8N�:�`��}F����p=ЕJ�p�n�AK-�rE�n~uk�sx��/�uϾJ����8uZ[��]{1<���k�5Qz�s�����CU���U��}\�v����4\\o����o�������� ���<-:�U����;�{�,m���i�\�>�:�Y��0���O��%N��T�B�٦?$�)�nL+��C��܊�i�KQ %��x��F�ͻ�?��g��:5�|N�E5�1 \Y���8�OAiuyݵ��L��,������՝V*�u�\����Ï=���Q��@�Q�h,��d������<�/�"( �'�X����-"W��fD][��@��^Z��S8k���vcejkN�q�Ȁ��,���2���A�X�󓈧�n�ĢN#�G�֭�j�0&y�/gql5��bWߴo��D��&�p��������v��[�� !�L`��GYt:Z���$/��``p��#H����b	�����z#��w*5,�>�s��߽�Op�U�cvn���W�;���S������o�y瞍�5|���Ɖ�	��J��6��֩��K��߼�-��Y�����]?��?�q><�f3�r��)w��<�1'0���4�f5���q�M�ƛ���غ���Ǳ�:�N������)�,�e�!���^�����F'�S�F<��8�ⴈ�3C]5��Yn�����.�uL�u ���aզ�SZ[XR��6#-ȧ�1W(�P*��3Hx�I��$���sȥ|�X�u��U8��TE��-�)����!#�p�n���r<��c�Ї��S�e�Їv+!�.;g�׭7!^SN@�!������/��?��[>p����߰���[5?}���{?�xrr�5O�����_�bLO��}��>,�ߘ�^RX�����D��̍�*�d�2˂���L"$���{>����G��#���kg�9K�7����#�[�A�R@��W�� �L0݂P*#�o�]XR��.d�n�
p*�k��=�8)ЩqL��hG�~Y��S�A�T;Uu�݉��r.X�9������x}ٕYTJY���	����ǝ���,$����X(�F��G�A$ҽ�CW� ��nDI��81=�%�:�[�P�L���QX<P����m'U��Wo^6�6���)F���5Cb�S�J�=1�����5i۵�H\���F�-���6���98�{�r":�}������7\��=�F�2)�
(Ӊ�\C���!�l�q�ǃ�cwE�
[�at(+\YX��d���ȭ��C�Uԓ�E�0���II�����ݐ��/*�SE�9��J��9Nn��t9����Q�ń��p]���@2��ь�z�\�?����(�
��lB[��P�|6'��K)�t��J��?����b㵩!PQV��o��,���LN���p��b��F����p��}�z�C����M�jU�a~��E�$ø8L�U�])�D$�?K�ݽ�!�����ϙ�!`���l��@��bS�.d�RǾ���r��1��^�MMCh������W��PXNI�a�S*W�8���4Z�A�\@��s&�x"���ɉ�դ�D�Q,���6"0�M$q�^C��l*V���!�V*�xe���zPφ���f�� ���J��!�5��0
�E��{E]����r)���y���s�v\t���A�R�m�Z6���
]��g��0�"�N"���&��k0��8�2i LG�BI]$k���9&�c�<���%�����H���|aU߫X��JsqeU6�1�q����0q��W�"8����~{���͵��Ok�t#]1���'�����L2��=�v
#�P*���ī�D�����2��Di���Dj_!6���GU��ܢ���66]�M<�'f�����(���O��n��Y�̈́�
�(C}q�s�p��QZ���9����5�5ņ`yyQSXNڸ?��9���Г�a��A�?���<��1�&��Z�f�(�r�6�ҜpB�X�`�,��X�=n�fU��t�|H��K�q�9g�9�|�2]�<~sǏ��4�P��&�m��L6�	�(�j!��h��K�6����j>�D� 
`b-���U�q�K�y��=��O�Tex�y�O�Rn	�D]}�##�/ӥ �z!���U%�!��2D��3pj���}�s��g���8�����q6Z�"r�'q�����<��gcnv�ꋸ��w��=�N�%/�	���W`���8p� >���p�}��Q)��4��M7]�w���18E��ƽ������ؿ���Mu��&z�����`��F��F��*n��9x�_�[��cf���f��S�U�R\����V�e�@�fp��V|F��04؋�~Kv'�����P]Cs�.�ӝ?rVc�I�P���^�h`S�+,,�\D�&p�Kӳ3����Q�@)�*x�=��s�#�}f��Jd����C4�@,ЅLl];q���q�Ç?�U��� ��C�F�B�R�hT/M��Il�Y̡�6]x�k_��7��-��ߢ!��/���g?��f8��}��\y�ex��'�o�ފ���hJ#�D0�/�7�\��z	�=	\q����׿
go��B��{�� ��{���b���J�&��f�<5�;��fWۈ�FIuK�/��g�E�A�Ad�;�y0D������榧���hM�QdW��H*�
��Z� �'@2B<�F�W��#�@�f	�FY�`��
ْ4L��IZWN�<�3���])t��#�A�XE<�_0��M(�nw0���R�j<�5����
��ӁFug�`U�FC���졾B���-���O鐤t�rY	 �^�NG��I�i�7~N����[���J�)y�8"��J6鈎dC�bZ!����o��P���?z�"�憀c^wL2V��ߞ��C�77:���خ�E��B�beM�Dx|�u=n�0�j�jU������}�)���h>��Z7gY���7�B��p��95 ��)�������(&�*��r��i���H0��	��lb\+�t�F��_ȷ����H�`���c��H'�I�j��me}� �,�u ��P +ĕ!�Qؼv��z��dQ�5�j�_�M��D�r����5�,���r���=�b�*��G�����A������}�~�4$v��Z�+�c䡛nAt�-NmBTo�T�3���޵�O^Q)�g(ײ�ȯ��D�H!!6�	)j6��>wZ�.���{�uR)�^g2,��vm鶢��=�z|f%�5�A���Z&��G����
ͺ�N۷o��m�����氼�,���0���.{�M��0j""�k�y-��d��
�n��ygSI=Cw]S"(���>i�+M�>�Fe����g����8i�z#h����Z��P�c91,�]��@k��A���;1��(��~�|~?�S%M��A�)N�lrM`���׈�SN��E�W�Jk��/V��Yl4-��h��f��+N��Y#Q�%�('���MSb!�F�uBM�}A6%L�f^�p&��HSO>�����gA�    IDAT�"���A�R	Q�<�pf0��k�b��;��*9���]Fuy	����+@�t!	�2��I���c�PD%��|����2��F��W�Tfʢ�ר�?W *-H����..������c�S*��b��!q�9�6��\`n�")¶���<K��Eb���J��㫫�(�I�����O��z��Q?�ӳӘ^��Z��P<�toc���đ�aAH������36	!�B��6��<�S�x�Ǿ�_>z�U�<��p����4ιd7�����q!����2���_��R��܋w��_����?������|�'h�\�Ą�eUE쳮��~�;q���n���?��?�Y8p�F��x��J�}S�����"��ny��ַ�1������r�@��R����i�:�٥	����
t�wޤ�R�}�`tl#��2����t�&���n�`gO`N.�+��3�p\���3�@����`H΁j��1M
r�&gg4)�B��HI��<�7��Rꮅ��63���0��A�݉At�GћŮ��q�7���?�MLΒ؏v;�L����࡮�{S`���Gem���/{����wny��������С�|�+oٲg�?��������y|��_é��ǰR(�Az��3��}oF�FMt_���ع}ox��a�7���"� �6v��k�B���� @���0�,��=��3%�C*��<,ĩ5�@6<K��%�F)�mӬ+���֛��mሉ.�x����!'��Q�o>oRF��i+�5�Qǎ-��>6�x4$����
*%&�$2eB"���(�!2�[)��a%�����rE�䊨4Zu�}&L�k�R^E+��9&%��r(b2��1��b��w qC!UGŤs�oM�������%�Q��r4Ŕ�F3Ǐb���&�e�nN>C��{c��"N�EK��Ԓ��.��֡��RC@��,�g<�\r�5�D����5!൐�P��͙{ D!X�7�K�����¢B�̡��f��󺒲So�(�}��+ҽ`�JdFW�g>gŴU�j|<+W�oU�q-̊O5�,��TE�������\��ϯ7l"\��'���סx,��*��L[E6���Ԫ�oQ#���I��F62r��F��"�!�}���#�m��Ǎ�-��CU��#킩�F������MK����o�gs���G�5��xY�q�z����1^a�{�5�|���΍�g�+��l8oy�A�4"�<��l�5g��fg�R"���R�6����5�,,i_�&#P6	ך�� =������J��=)S�#7�QԞF�_v�ɻl���E�*�u��.�F�^�YZz}z��3�=�Q`�xoǗ�4�_�u)޹L	̉̚G�"�U��{��9~=�/�;)#ٵ5��e��|��s"��1��0�="�^�&O�/��X�aɻ\�jl�ia��Vg�YG	ȥJ�٬l�I7���'�e�{��B�B�5z�8���eMAM�l(�P�E��f�mk�>멚=��[�xI�I!�@�H���|�糺6�PTS��!���(�Kj���A]������'v��I�U�l�k.w��Mx���%n�p ��DN���׉����ԡIA|����8FR!�:��=� ���&���kNg2�^�s�j[FG�m���r1�L,��߇`���C��K(.-�������2��η*��P3ky��K�<B3	��+�H��XE_*&mƥ矋K/8O�Vav'}��e}R;�,1�L4�zC�n�_>+<#8=$�W����Qqzu㴭q鳯�஝�DX���ajn+���n��?͆���~�AQ�#о�3%E�#���щe|��_���h��h7�R>B�T�q�E���s\��˱������K��GnC)[@��1���ߌ}�����8=�O��%|��w�U���lƫ(�06ڇw��x�+n�)��s|�C��C=��Z��pW����0S��k+���,^��}x�_�	�]C�-,�m��`���8|�����Ѫ�Ź�"6Y� 	c��Ai	��ϯ
����Z��Q�%�.�-�z�l;����<��aR��QR�X�xRzR1W�VU�؄�E��w&����0�ܐ�B�^'�'�ƹsm���ۦ��CW��]��M��7�[��⋟�>��ocn�,�^�|� '5Y�p
O��3q�D��N��ja����_�����+����4����o�}�Y���HZ���	��f��̯�D�	���C
�U�HHH`�DӀ���ɎG�����64x�WM�W3AkN����>��ǗN!�;�Z����<���:I�g
.�34�!N�]q�]��_�XR��n�RN��N�I~?�����}Q F�Bک���}�N���W��d��[��eU#b�6�DW�###�?����!6�H/_z�7��ۏѱmBh(Z���P'��*�d�6�d�P���	iZը9�$LyOE�_�2��|��Fk��b�b	��:���G]0Y��f'�k�ߚ�'��ϊt�D�Xs<�]O�5�s1�
��!�������E�����I�Qf�_�e
Qr�1|�U��G� �8���D����RO�z���ib��
��i(�-�8z븷^C`�]_o���gZQ!�xt6$��R	
�q�^o���� yӤ��ζ�-�9������c����IRb��u@h��1g���<���fSs#�E��9;�h�6�F��^�Qq����t.�������9b���ʐ�����;S#a�՞Y��_)�<��  z�����(L�4k?pfq��,x^�����k��8pr�5�	{��$��n�p}y�6�l(��������1�t2�7_��rH��*ڣw�İ���0� ^G~��L��K���/��x��,��8�>,�Mxe����Х�&O���R�fM�K�鵜~Fn>	����u��O�	�]��]�M���"6�N����֦=�Ds��=7�8=	�&�!���h,([�b���oj4���p���hx�hB��/i-�Q��"�I^c�lKf.K^"��������%d�o#�A�I������!N��ӅǛR�P z���q?!�E�<!!P��"���֧�^�-g���UA�7�T�O�$�Sz���0x�)����iZhV�NE1�	a�G�x�����	��fW��<66&�%iiL���35D}y��5�ۍ8�r	}�4­���V���|��+[�H�X
��"��2�i5M��M3UQ�ɸ���x=�����8ꋫ���*U����n�
�r���\�h����?6���P0��b�TBm\����=:�R�)n{�P������!�9s�MheY�j*@`p��G5�4C� � �m;�N�㓟�:NN3�+%� �8�::Lj\[���Ļ��/p�uWb~~����/j2˽�����7��q�9{p��8>v�W��o� �]���V�}�^�����o�K�A��G������2�E���Xʄ���i�`���Tl.��5�����W�fl�1�م�ȗVI�P�����tȵ��Pa�W0�����cfG�-w��E0�C��l��,c�ܲ1Q��3O!��̀B� @ОMw����c]+ �K��X�f/Q����/3��ų��ҙ�s���q���� \<.��O�Pw��z]�s�h?�C�ڎ��.��|��o��wރ�K�9"����^�X�y���sA��k�������]��7�n߿^�s���������9�}�疛�B�!���|��V�1M�ָ���ؐ�OOx�xk먣\aQ�q���c�F�-�9kN"C� ��TB�^j��w=��O�"�Afp	Ry@��;�G.!s&	ț�I(+�r��Q������>=��o�(SAZ��Ŗ<�u�Y����Hr�Ѹvqnuژ�"(di��D(�A$f�-�zS3�ӭ�J��kD��(�VsH$�زu�>���,�[��3�5�,R-\�K^9�_���)�U�C{$�f���oX��{ra��B?�h��DŇ{X�Qm��H|��S�f�8��*�wϴG��k��A�?�l@�t��v��[���}���#�k���
��)��Q��]C�"ːP[#te�\�j��x��ZnT�!�^(�\s���G�QQ�Ę���%L��ZL������C
�I	P��cC�QsDGp\e���YA�5B2�����Y1&��RTD7�*�q�Ձ��k.A�T7)�M"�H��A8��:|�Fsה߇��Ffl��{?�H����e�!�Gi��Ī��U��P*��<k�"�Gs��L�|3���ǻf,��H�Mז�9�u�ֽǵ��s�v.�1�u#:��'���s��@���0J��
�����=19E���1���r�h0M;�C��k%��M!x��l�{��1i��Od��h��Q��i�t��ަ/�ӏ��?�R�L�f�VH �)Áhe�=�k�G�XP���_]c�B�BIk=�U��T��2Р&�j� �f���	n�jͿ�]{�Y@s_g�gSNF�i�v.�dkT��!X��꒛�oը�����11�G�}c����<`{I��N妆��F�snM�����5~_H9l� �w6BܜI��G�l*f�䛨�׍Y(�Je'A�h;�L+��e�ד�ܴFD�i�D��$�sj�T͛{�=SrY2Z%�%�\�����0�c��cUWq��?�]��&|B����!=7,��IJ!�B��}��0��������e!�[մ�;�S''�L��-2q�4b��k(�f�C|�n1�T�}<KHɡ�+]�H��dnJ�(;����#e�W�*Rn��k�iA:I��&��&|j��
{��j���YWc���X\]Q��T���y��s��>� ��7������Cz�*�8�I������sp��4>��/c�ԂB�X��~��`Ӈfv	g����o�7<SӋ���/�C�M�r�w�û��v\��+057�}�'p�w�&.jʹ��o�$���eϸ��߷b۶m��]��m��y� ��E�d���MRe
��]Zpj�n7Pɯ�E/�o�����]Ø^�@��G�'����8�(��<�jhZ��!J_200�Ɠ�m�VC>��C=�WFKem�Z�������(G��B�$z�	������d�jo�M{q������M���1��s����zE�
#E-" ���H16G��j4����@2ԧP�mCgcz<��o�~tϣh��ݛA���3�uS�~� ^<&�zN�Z�T\|���}൯��_=<���o4��>�[���;p���_���"���w�s�/>w72a+4�0:��a�6B2Lc�p c��܀9�c�?U����ӨV(��
!*���-��bxh�2��3?@�A��=�S
䍍p���7/����"P9D��p�g��
-Y�J� ����ƌ1�Z�l@\RV��ɫ��\��e8޹�Hؤ�@4��z+�ZӍq���M���Q�ǲ�b�̓��Y"�C4	��m��%|3���_.*N��f�E3���P,6���
�5�D����,!�q���:1��O�r�d�*��2|j��U��8r
0�łS<��`�B%�P
���C�MB�ᖛp�7�!89?����1�@�A�
)+��������^衟��U�+���;�km��si��0�o�w��%��MpD'q���Fz�**91p�g�soݸ�ڞ)ϓ���G������~kt����3ar�&>�hi��hx�,~?:%y�f3�˂X�I�(&�x�]�[{D�y��ɶ���~p��k���*y�(X�����!��g�='Q�::��B�bW����9|m�ł�C�u�h�����2��_�v�G�ژ*�B��ܴ�U����O�x��+e�I,:������y��C6��n�j4��lI�cS��Tq��!����ծ���9��[�B�~��K(�֥�j�_F�b#/�6�_�Q��\��a�lz]�=�5K�w�	��C� ��ߟ�Xd�z#�MUL�g���F=/�
�r��`p�����{��G�J�'���ߗ�rYr�@!�lD�sf2'�/���5lj�Dў�C^S#3���y�{k��FԪi�4�)���r�2l�.|O�sm�"l�,4l�����`Q�I�Lī���XT��i1�=�}��
8�#�/|�3�TA!��>��D�R�Z�`"�x���S�p�~��/�;Gp�=?���|�9�v����A����{�.��ӭ+���������έ�068�gg��i��q�����b�x��f�6�x�#��/כ&=��ɶ�%�qr�X3���¿��pfp�k�l��ISWBG$�oH��6�� �1<oXtrRV���c��ʫ���o|��&l&��<N�:���)�i�h0x��J9��عm���r���qhl�(C#{�����֏��Բ&����n��}m	{�ڊ��w��k.���
>��O�3_�2u�u�9c�W�<�:��E|�_��~x�&�����l�X�{�3�go�#�ڹ�����������P�uЪw$�U��I�M�T�8#��VE-���t���{�܉��I䊫@��|;����q|�8��5�y�h����appH{(����5T�E��`����t%P��P,��Ч{A�B8!��D�Y��C�j�z�:Y���H/�hr܇�3�k�\���"��@�����˟QmV�`W�j3�x���?��1�ret���OmEo|��F����w?����X��Ȇ�I��&��5Ά���7�Z	M^��j�կ���7��K��ߢ!`R�G���wN�/�����ܳ�e���(
�H���@�B�0�o�Lrƴ]-B��1��u����K�����S)�N�.��p��?{��𥟢܈�wlB���n�>"ТΚؕ`�_���_eH�G����.n��9���67���U��p9.B�t�n��F���]��F�<�;|a���������DBE1�c:������UW�=8z��Pc�c�C�W�J0��υ�Idl�j��x�L퇄T�Z��3��"R�҉��g�'1w�J��4��O�S���z���������W���T�h�78��'�M�i-�H 7��x�M�SCptrJ����CV(��B�C��x�펏�9
��c&:j�悑�Whڵ�{����1����a�d6�W��Z��v����Ԭ9�o��e�xv0�um�z]�P�
!�lQ�~��y�+{-V��pvBf:�z��^ʮ�&t�?\��]PD�e�	�HN�������S'B���2J��D�`gsO���$.�OAJ�מ�.�n��@d��� ��2�hs�����޽�i�P�`�jC����5�6��s��"Ͼ�M�4E�TN�M�6�'����(ɷ��b��"Ŏ��cff$� 1�	�י��deo8*S$�\G��sW�Ll.F].��k��>q�_ž�`�[��� �y�šw��|�t�=�ۃ�,��΀���Q����wUlcvp��akyX�&���P��)�I6$n��d�{�s�5s����&E��<�)L��v=w6��v�=���]�&1<m��D�,�5��u���ߢ��k�'f�e����/�f�(-���B�%6֜3���k�}Vw�5��� ���F��j��UыXs�?�й��E9�����}�4lL�h�(���i#Ѯ�S��MϺ/��*�EЪ5�|��v;��V�ަe4�>��b�^6is�Wq��8��fП����
���e���8]\YC�T��j&_3���#���N�.�4��%��E���H�MH�ʺIf�cP[4��Y��Q�X2�PH}��ղlO/{ڕx�o�Y�����,N�<���E"�"�fp+����AlU�����b�
n�u����C��/���&�6�Gf:Q��A�RG���Y�l����w�W]�ӓ3��G?�;���,u�.��3��y�[��Po61��G6_��BJs�h��� ≈�ώ�[�l-/�`qqUY!3��8q�R�]А����Y�FK�N�Å��X    IDAT��)\x��xӟ�	.}�EȕV����B=�l3���"f�f��]��ڂj^7NR؈r�fn���
����{咔N��,S�M*k�9 �)�F-�T/c�����x������7�8'=������5�v��)�����P�D�I�߯�c��M�?����3L��t��Ewl��1�$�!��7��1>��;Q�s���:6Ɣ�NZ���Yˎ��zi��B��/��}��×���##˛���ϿՄ���'>�����C6<28466b]��]~����XR	�%7,�]�'�C_�Z���۷��3�R0X8la����Ձ�:�;��(r� �#�ѕG��5:�Xa@�l�����fm��<D�a�DLC�x�P,�.�Rm�X�OvE�@D�Բ�QAb�'ȴBR����&�Q`U�
��X>�n��T����Һ�O�z�ʂ�,5.��P9g�����A/���%�isN/��	f<N������J�2uQ���'j	�OM`qr
��Y�U� �UC��$L{�ژ��Y�	��$5�Q��x(q�x�4B�"�3�5q�-/�57� �P'�gQ`:��.g��P;oZ��Fq�Įh�^u�D#�u��w����eC���Zw�q\h�ʎ��5^1m�Β�̽�k.HѰ�`�=[�&n���k(D�Y�Ys�>�I������5�ހ�Wn&�@�\^�ؽ�+������oI���H�Dj��@�u��U�(i 6^;��a�5��ă�E�����c����!�*�L=l��k�4�5��W�[A�A��6G�mW�{�'��O���E��K*F�V�v�y��>��������֐'uii����>����$ȡw?Ci��B�\�):���т��8)��4Q2@��*���,���OBZ�]������]�!G5���lE��q~�Ҙ�n��D�A4E��~�sS+�Ul"F�6�� �GZ���yϊ�{�5�^�Pj�j�L\8?p����`h�c�u���`sX�ЕXٹQ���kD��s�!��5ql"�;���	�i���o3 �k(��l�)�6*���sx�	�,k����p�V��I��D���ɣ�i�H^q�ϼ�97"�k'�_0��x ���7p�� 
�|y�>�l����MS��@��t�b�PXB��&Ͼ�U/���;�`]�>��~��89qچ��6r�sl61<�/��d,.
R�QG1_���6��������TWZ�2Ӯ�8p��xR�Q�hBAmN]�Ea��WMPt��/��M|�����2'q�:�{�rP�X�MM�����7��q�UWI5~�8�8�3����_�t��s3r�ZZZZ���À��.�������OM-�iaLM$���=�b`dx�)����1<~�$�u6�Y�p�0��T����?������1>~���K����#�-��c��~��;�/�w��"�� d�J�!>���;+���9��lE�ՆD��h��G,s���#�L��"�k�>�{��)��▗݌��4f�e7:���b~�˳X�-�P�"�=8D�O�=}���
�YX�C��G*���c�A��e�PO!�*uh�)��Vkב/Pbv�X�;�6L�7�4�q�4'h�9,�������Q(��'|&�{�ϡɃ�\����Q�E�/�x'��� 2�a�$��'�����;~���a4;q�~Bq�Cq�yt#=0Q�e0J��|t�[[@3;���W���?{ݫ?|�Xz�7m6��ߪ!8t�P������}�ɿ����C]\N?����)��Us@`�h�qs��q%�X:����i��|��/��z\xΙ���Y��I^ԁV�<qx����V(��B�w�pi���4VG�����\%���D�a����W�h���ڍHG����D��+�U���ud�z�+���=Nhˢ�e~�D�<7����&�0Z�-r�թlH8�0.7]�aԘ�hMJ�u"W+��� ׯS�C���uJ��W'��5Ug�ڕ�#I�)�W�6u�4�������g��'�^+jܨ���lY,ڤ��H�8��W�i��h�D���K�c?ο�\���Jc�TPCP+�D�b=���&pm�Hu�$�����ڨ�c���w�l#���:
oc��^H��?�^���@�7�V�xV��C�7�^C#�չ%yk�E��x��I։^t<��2y/�-��8{H�7�)�
_6V|����ikD�]�K���n6庡p�FU�!7�Q�!s&��i�H�4 j'�<t�gs����h���i<XXQH-�K�7���5���<]��(xMIXظ�3��#��o�缆`ݥ��2�����,G;No�Y��⏅��*%�	'b��[�[G�Yo��#�S"VܟxI�̺�3N��$JL�5��y�����6��haͲ5F�Tf��{ͨ�25�?k��{.�:�h�	=L���$��9��^�����,�-��U��֑7Y�A��P��B���Eٳ����]Zb�B��s����Ntnm��$�vS_�}pQ���}���#�{���7rqυ�<3��� �"�u�M���l�d�#���&�uq���$7�FǬ}7��o<���_S&�i���.�Lg���D����"�%�U���::��9���D�WKuD���(�_^�px�K�������S�Gp��8~��_bfv��V0�[�Hė7���\��dZ�6FFƴW�&��v�K��?ý���r�x� ���لќ^6B"��qN��%��+m4I�ؤČ7����I�H�4JEݟ��^���	����Us��'���&N��p�%�+E9jy�F�V��ر��{��mCW"��+�P�g�HB�}�c��C�����!<��(jM������hU[��r��3��\|�98t�(���o�{��)��i�0:փw����� �XP4�em3��go��)ڕ7A�\n�6��^�Ǧ�����_���p�ؓx��������N�fO`|������[R0Y+�B �ku����j�H5˭���Ė�D�!��p��癮W�V hďr��烩��zY�N]��pD@�Q����3��a4�S�iM+��NQ6����AE�t2�����!� J#�A"8����ķ��{೟���ϡ�g&]�l�K0��A�9,���8�a��h��@%����k^y�{��5���ӷt�n.��?�VA��������>��?R��hO:&��E�)��%�$mn��f"��!z���Q�ʋ7��^���A�������@�d�r�سX����r��'�����ca���?�p�K�H4��/*��f>�:*5�����핏w�VD�ZQ�?�Zi�ɲ�Z㘨�R�CruX���m�.yv�^�(!'� ��Q�M��%ٶ��h!�#��!Uǉd-$lÂ��qW��cꞐg9߰�k!���v�qZY�#�K�
H�:�VA�d�;�VBB��z]�J��RO4�XY^�\�X@imY�!&�qB��\3Q�j��B�I�`�/�4h��O��Ʉ(����������ٗ^�P:�|�E��������������F����^qh(��r�O���r�q%b�r ~-�U_�(�C�1w�Ch�{&��z�����_���ӏg�jE�F���'7�\�d���,�:�4kAZ�I��(@�f������ӛ�y� �x*e�H�:�(q�k�l:oiצ�w��-����%׻��.,L7�q���<;�U�g��y�F#���
yM�w��umx�{t#(j �wR��h<��օC{]�Ͽ�|?�"�~�2��B�H�$�t>�94�s� ��G�s��zݼ��5�E�n��������w�^M�����f��~%s�jk�\�,�����|x}ĹvT+6C\7֜l�ܛ>��:o��/�ݠg��߮�������L"<3 �V�MC�3W��#M����F�V�ю��������gD%�v@�{�k u�9�����^6�T/{��my՜�ꔖ��PL7=����D�8I���B��Y2�M������Ĭ�s/��	�f�j{�7�6���刖�����;��('�ԕ�Ѧx��C
e�Q��4vu��0q�&&O�Yͮ![���{��,g���+t�Ju�u��b���j���^����������#XY+ȍ+�[(�F��$�̲�âʹ:�DDSh�?�
�2p�sGc���OJ�e��fr�$Q~*Ӎ[o����$����"|�A���h�qz��� hçٝ�|�lv�2���s�Į�1��+��B6��P*�F�|0�L_=>���?��_>r��g����.�m��:����½x�{ށ�.>O>�;�?��^�L/�U/cx�K����f�a���@.�G_߀	l4Y��M�SdN'����������V�����H0SY �AZY�}��}�x>����o�ڪ�� ��{1�Zx�O=���,����2��
�^q
�AO/������U��,���۷��;�����v�/�6m�*z%�� :���>�P�}Saf����-�Mp�г��E�n�&j�*U��Y��$��u�Eӂ��v��Q_qZ�b�?̽g��gy&zWN�]�{r�(��HH�%��� X����&{���k�>���$�	�P�@%P������*�:羟��nq�?���K�LwW�����p�d;�5�1䓣H`�}�Ѫ����?��N�T?�U�(i���Ŏ-e����a�$y�ct�˨�W��o����o���7��'|�}�o?|ǣO�}�`494�n*�lf1r�U��Ӥ�4��`AUD�@�e��A*]�6�cm>�M�y\x�.��c#�.
ˋ"ʱz]'$�E��/ދ��|
M�!�F��E���ÈwS�$�ԆギS��^��[��֎�b�T��'۟�:�6�6�3����:�M��]?�TBB h�+��J'X�#���+�@�@E��T;Y�$[�)i�7Zm,���i-��`0T����"�t��^�dW��%�Y5gEJ��I$�[u�.i�m7����m�l�T,�U*`��a�� I��"	St�Pi��S��a���#�!bɭM��ĦMF�Z�f�@|��ظ}3�c\�J�Z�gQ4� &���f�q~��7���U��]���Y��3!P�8���^�f�A���x0�P@��!�\�����r���ѫ����(�
��ʁ��U�!�,pS\�1��LV�A
�!K���ԉR��i_�|��g�≉W��b &�$&����Zf�e�zUyv:z��A�Թ
~��.I��+�ϫ�
�B%�]�� ��������O�WH���`Y�d����ҿ"g��!�"�qO��l%�������%�=��I�k��m����d[$Yk{wY0�^��8A�}��k��x���U6l��IL\e(U��3e���g 跃���S):3H3�W�}.21��]��X"ʮ��>^�7�k8���N,)_I�W�0��Q>c	���X\Y�SH��hT�f�';����P��S�����9	\r�I����4��{Y��O�#^�W��h�9c�.��Ʉ�)����˻��C%�D{�.���!ut�FF�i�N��A
d_�#v[��422$%����<�KD=�6�P�Er�ܧ8\��D.�Z�%A���D��}({	}�:��s��>*����u�I%%���/��v���(�Lg�׾Di\ߓ��r���C�R�!7��V���j�)��҃�[R�4��r���Y\8H��|�.�LT�ok�c%������⋅l����ާ�����⢠R,���h�[u�����-04�~��6n؀5CcXZX|gddT��<��>�~�i|�O>��o�8�t��v&�%�yƉ��W,!xf�^\y�-���0sl�Z	������x��O�m���w��x`��յz�D̺[��'��]�v	�x���yz�x���vH&�VN�*�/21	߷G�Gg�<�_>�KL�N�ވK��Vt��~�iD�4�+c~�<�Yy�p�e\�dp8?,H�!r�)��ϊ��n|B��f�"��,�X����"��Q�hR���@+֑��`yV��9�|� �bJ(�������?��L<��ު�1�K�8��Y��s��3��"X�_���HG'Шf��c�p���a��004�V7���%i�F39Ź�S١�r�	:�Z�v(3K��ť?���}�����o\[���Uu��o�����;�C���Z���a5���� X�Yx3�A��x>mV����q���'�02�ӏۂ��6��u�X?�G�ۖK.7�j��r����(b}Y�v�^�p˃ȏn���0_�`viI�ch&�K�ə�/JlV��0�V�TZ�Ɛf��O�A�<�XJ-�B��G�s��C2��9��h��*`�NSMH�tti��lT0B���!%�d����m��F��"�d��)Qz<@-!�,v�u@ǩ�gɈI0�niU���]���@�C6``s)�K�}|a~Q��H����$�QbXIv,�I���j�*�i.��Z��X���12>�u[7axb-"�A���f�rV�ظ5:1G#X�VQU�A���Pywؓ�U��W��2����WND�@ǃD>'V56A�ȃ2'*Pg�E�V���b2s���0�F�P��ʡA����i�������P�Z��F�l����dV��bm뉶*�7nT��	��CG{A��_)NY#Y�*�8Y�8,� i,�:��$�d�m1X��/��%3���J����}�1y0f��t�LM=~��\=N�+J;�k��W:|L�ga�v���ú�Wt�6��$	�"�h��X�E��}+�ւ&�L[�$,-�'TB�0U�١��۪��1�.���m�$�����=�:�C�6��B`')jJ:��J*ufԂf%Z�Xݿa�eT�mUb��WKx�L�|=y�C�h �[�h���(;`-9F�9�9	������?�n�u��Q-'H�z��֌%Nt&.��P+��a��>�e��DN��xģ�P�:���dI��=V'`~�R�	][%�A�X��"H0���t��6��BǄ-�-�^'s� �S2d�� � $({I9"�H���A5�G�Um=x�HOJ�KD�����]r��Vj�Zn"�j!�*���<�dc��)~i/��22��C�*4HF�~ m3��t)"�%`	�'F|�wV%�V�I(X*K&�{cW<�������s|A����K�D��N���_�C��R���x:���k��g0;9���Y�c)����Le0�f��u������ظe=i�X.-#։btp��mB��t���G6�3]�DϾ�2~��Ø[*"Jiv�٥aW�N�ZB�Nė���8�����������]wޏ��ڵ
6o�g?�)\���cfn߿�Z�p�-HQ!G�TS��n��p����?��T�~��1����3��5Go�WG�l2�s1?��E~dhX�&F�'I*}l��t�p�wa��2��e��P�pt�0f�g��GC��|#�#�naqs���Q�r�I'a�ĸfC&C_��U��%TkE%�V�;�eg@�DW11|�8�L���w���j�� E&Jo-�&"C[7��4�b���E1�_���u(.&�����Ov��� ��!�@��E�!��G�:&�>�F����P/�VhV�Ԑ�T���C��o{ەgo^~U�@x�J�!��7o���{�+���!��4jى�&�hKK��6�X���-�}���Kyͮ`)�Hù^w�)x���-�J� (.�M�|v^�#㛰f�Z�yߋ��ǿ����Գ��B��}�`~��f���I����fU}2djQ���d�����:�Z�:��������]!N<%�)H��!#S��щ�R��F&�QFM�XF��ly����C��P��7�٫����aupK*�/
LǿW���B��*-�gVe����'�1���@�UCU�Mk]�E<8[M��寰0;��aif�n�&F��O�ը`z�(ff��ӬchxP��n�    IDATO�#k�
��Rc���L���mܤ���m) ϒ��t���O�1[(`��H�d���*�VUm�0����,,^P�<���� c�è]nD!P�D�p��e��'�	�*�l�20U0�.�%g�#�ip-o��O��c�W��+��^5ڱ�ڸ,y��W�4[IRԪH�Z�K�G�dD��`ǎ����)���˚g�jz����|�	-�
�;����eqς�:w#S} �z[.rm���p����J�y��6p��g����`s�sLF��<�����p�=�Qu�1�*ϫ�<�n~ߠ$��F�+}-!pO��f�@�Xz�����Q7��T�P<�B�a��X�H[��9f�E�VIw�C�#u荫mI��U��K%,����h(!�F%9NШ�	������)Bx�W�=�C��x)JH1غ-2����Y���` �	ǐ��8�˦�L	e��b�%@����N0�1Q�k��!���"ޠgI�4�G�u��D\�o�ާ��^X�@Ò��uq��(W���� r�w�������&�O�_t��.���D� gw��J!�aW�L�k�8��`������y���~/
�y�3��{X�+�8DIT
U�����/�[��H�����,��{~�'ۍ6�!�1�>� �sM�St�6ވ��B�G�x\VT��}&�ɠ^("� ,@ӿɡ)G��Ɍ�M F�vX���I�A���U��(��/��q��N�(�t�>�Q�����b�Qo�:H�h�/Y�!���ۮ5��pl���ڢ�w�zM	��M�Q�177�r��3y��z��%�V&ׇd6������Hf�]Q�T���|L���2��u�������N��߾s��b��N����7�?����.ž���+��o�]�G��s��-OO�1�_~9���/"�N�����?��GZQ$�݉��Y�X��d͋g�Ը�G:�B:�����e�ٺ�9'6l�#�&��N܆J����^��C�P��U	�46<�n�$�ݻӳ�8��m�&���s:C�\U2*�(Pm�Q�WPGu�yF��A��{�p�$�-.�ס��{� �K�J$�8�H�|�Yu
bt�xMӹ�R�Hv��@����_���?��ۃV#���J��u���������ܻ���A�e<˪�-f��O]v�y���~�{��)��'7<����}���>��?�Кlbhm��버Ig;(�x ��f��,M�}Œʸ�����78a�&\��ႳOF6��D�%b��b`���#7��?}w��Wh��8i�9��d��b�l}�Iժɥy��a���T:�5k�m�.M�ծkä	����6 �33�869�V?E�_2���_���Ϛ�@:��t��N�rQU!�7E�lp�j�``U,�0=5��%Sr���UMƑVO�A���#j�S$T�J�.��� 8��$v����#���� ��c�l�j�Ę��cX\�C�/���~\x޹Ȧ�4�������C�c�v���J����Q�X�N�0�R[��+���� ��T\���RE���zK���Sh�#��e@�s�7>�n���A��{vH�N'U~9���S��4΋��t��Ѫg
�X��J�Ϊi��靗T ������K\v���E�D���)禒����52$��X� ë��-)����A�o~R&מU��R�{q~���1`�r.��:�[.T��J�U�$�P	�ɇ���*�c�Ju:���1������*�P!�L%S��~t���\�=]u�"�� �&V����k���6s�2��x���=�����.U+���a�@��-�@�C�9	k��C�^�q}*!�q!���G�&���}���dӒX��g��cɹb�K���u�QV%��� �Sg��iaN��#r����T��^W$�����>ל_��j��\�xe܋.L0�}n����sHVXmΐ�DIPi�3IJ����� q$�������}�zw2��"�I&���x�K�?�ݶ�����{	��u�+(Q�@�a{�';��j�L?�.�T"�Ԩ��F�d�?�5B-��ٜ�[��,q"j�-b�C.rnP
~���W�yĽ�R�h�k���4�3^D`�V<�֙��a�)�*	/�ϣT�#�j�/ZE{�0N�6�����E����?��ؿ�"?;�J�d�!����XP�k���ɣzFJ�#�7�<�ѤCp��R�cFMь�����h���1>kq����_Y8c���м���ݯ�o���ޠ{o ��~O�wmo��^mO�f֦����S*���!%B�I2ܴ�#�,6lڨ���[Z\����gg���Qr2��[S�Z�8�c�0�t�h,Ma�v�K_��8�S���}���;p���`�Ф
7;O>���'p�_�CS���o�u7ߌ�i�H�(jRB4�����n|��G�`w�q/���������U�H�T?�ev�X�`Aa��K/!A��중��B�Y�Q$G2���my���s�߀����+�<�D6�BeY{τ�1�|ڰv�:��sxz�3R��:�8��y&֭���("�6*�"*墒�B��
?;A7�����h�e�A����kD�1��T�艔ؼa�M��@6�D�3�d��l"�Lz �� F��!���n�w��a<��!,OV��ax`\�ކ-[�;�{b�n��x�hw�B��5�k��v7�����Ld�?���Kް�_/8�D3�x�_��Cp�CO��?���x�
�Ǔ�<�}L�$1<YG	��,S�T�@�1g����t�lС6�t"�f��l<�Mk����5��01�-�cӆuF�f_����x��$��`z���%��EI�Ku,,,�&Hh��e�sX�~�>�����˪Z���41r}����fu �_*,[��JK����k�r� �M	A� 1��*�k��^o`~i�bY�!�̱"6?G3��ԼQ�&�>Ӝ(=�j���2��{ qqA����vpG���KD��s��k����@���tǎQ�D��SN9	�� ]���R>r� ^z�E�3)��X�����0�Ŀ�ZS��)/��\�R��H�Y5�h��M��C8��S12�/�?��}
�H;N:#�kT-�k4�t�\�+�a
������,��@�**?�u����*���r��Ai�o)9� =�!�͆���F�4�>%J
���ǟ��Mp�:#��ì�		��� �ڨ�a2�RvP<i�����K��Uh��]XR��=V$I��6�4's��]��MS��rn(����)�y~_���
��ڔU��ҧ���A��%�����	�m��)����$F�5x����\�`T5�*v�C��a�F%2B�	��+�eWL:�!Q��ρa4֦�tq�?���9�Q�D)�Tp�@�{r镠^���H>3=�|W��e.�#�C%��)	��1!=��߃'||*�1+��䌴I�a<��<%�LQ�9tr�X�@Ġ�k��� ɫ��g� ���p�L��$'�y�Ġ��y����]?���]Ak�q�����ο^L�������;wY���:.4{�9�`���H�v�+����y7�� <U�[����Y
v�	�Q'@�� ��1�q� S�=v���IRn.����*�i��0���5����GN^�P5b��/7m�� �	qal_�{3 �4*M��)�P��?��;q���C�p߬�2)�!�Y���ʥ�� ���9΄�I*�m��=�m��:B��������/�����ǑLF3�]/JrJZY�7� �����G:�L�U���H�H�n����H����%�j[��fEE�NiI^<���$���}��Q����v;���A]��L��E�	r��I��v%+�0��%����Y<�"��i�}����~'���<���яq�]���\Rc������i�����c�q�Oo��tf���0������z���.�����0<2�;������'� N)��a�j��hxǮqWL%@��������j����m�������sN���q)N:}&�b��Q�/cny��E�9G��hM����
3�&g�077#��uc�رy+N9�De��*WQ�_��d�X�����͝x���ϭ@%��(V	s�-���%�ɣ2	JP%�A*�Vw ��!�"�C2я�����O���'17Y�Q�F�~�V�;x'�~*>����8���F��އ��\�lc�d2�1����������ч�i��g�z����޾�?2t�O���o����ȯ���G�鲚�E\ʎ-�����%I"Au�	��ϙ����L	"v�Y)�۬�U�a ��5i��S�hxd��a�y�͎�A�:�nLM/c~���h��9�<x�4�����e>2ڏD������r2�x�Ǵ�1�E��Ĥ�?�ܧ$�M����翉͖d`�Z�N����l�3�-������/?���1�8H����?��8�^ͤ�W|�j�np|_�Kx��X_�b��q�����
��r9mf�cb�HF09yT-��۷b��b��;�#(��739���퓓#[��_f�� �I���`� '~����>��s&6�T��2\x�8rl7��s�/��u�	ظy;��(�(#k$h?p���o5\��h�-�u8�W#��CWs
I�%R�d�I�$V�Z��(I�ZwafG����LU�N�C#j���1WQ�'(��{�U���\�ܦ�է�ɯ[��h+��*=~���åX���d�B����N��\�ۧ�A���#����}�!*:n�������a��X�̯���{&$��$x���מ�'J5������<�}���ח��z���<a�h	�(\aŏj,$3��*�̩��ĞR��\
�F�� aW��J�+������U�eZ`�O��+I^u=�����۵ԙ	��ꍦy�����`��,�x,<���v7���4WԜ|\8����΁�O�=I�3 �?7 ϒz�	qp�� ���o�T���1.*E[K+u)�L{��ɮƤ��cV0����4,��ɞ_�Uۙ���!�����e�d2���F��U�1��r���v"'+�%n^&[ܟm^Ɠ��1һ%ά��9�sV�3����B�FC/;�b��Jؽ�z"����Ɖ2�u{�(2)�|�E�̟bA.���"
�%J�O_^�G�R%�IKZ���I���T�Z�#Y�jꀼF��%�"�6�,�q��_�S���};�ڹT�*��#��� ��L`,���3�+�f�(Tbm�I2��{�7���p��7�W]�F��X�����Dt��	M�����3�����w�EV�e��T\��V)p�|~��5����N�U�q[������Т1UgBp\)�0VI�����zC	�c��1!z�oj��3���״\D���R��A�F	�{6>���c��x�ɽ��w���w�+NB�T��m��/���<�����݄o}�����׃F&:�zTK��?�ןƚ�	�����������O��)ˠK�B�T0��5	��r���ю��,[$�f�V	�0�i��B���]��P�/���}x��X(̫�G(��Р���MU|!����G��bzr�REJM'n;g�x����&�d*ړk����j�����[@8;���L8�:#�'�����^��],���/u��u$b	��Y8N!˂�ԅ�*�6<��r�?K#�Nڶg�:�n?��ϱ��W��&6m�5�߆k��S��H'�2�l
ȍ���_�~�غ}7]sC!�h~���^������y����������w�c�Hv�:�d$9�Ĕ��"m���!0�w4��&�lXD1�sE4d8A�gL�l�XE�/�A�@_�p��@���H��0��(��8vtŒ�|xܔ�V�'	�mg���HM��z�V]r\������f�dΖI*��-���f�΍X���!��̉ō[Akh���O�*Y����4e���(f$VظQ21��� 	c�fR7�h�΢o��4=@�B^� A�a�M�AFh�b���km�Ŗ���ЮK�I�*!��I�p��S�X��5�v[8U,B�n�!�`��R�(0�N��d�7���p湯�e��Nt�	�s߃x���&�^�V+�J�/�a`���W�}sZ�y"�A�W?�a�P�{�j�.J��*Wܬ���7nrzr0�|?�dp�;��+!����|���\��J��p�e���7[�H�1�ܞ4���A_%@L�i��#UQ����5g}c�k�q*P�p��%e� �piEwY�8���0Ms�_�L#�ǫ���������_��ą'�J��3`�ݡ�}dW��.�^�[�QB!�0,vR8��jo��2�VמI�3�Ù		֞Lrl��?vlR��d���!��l�m�r�)y"&�@�:?r9�v���)M�!�������1'4��F�5ּ>�T�lhPl�`��� 1&�GvA�~�W�y��{�|���w�<�Q���0���m�B�8N�x]�+�8����тe8I�v�al�`�'3��upb��R6?3���)�rY�'(J�h����r��{���CI��RQ�[�A[�R��s�X�kTp ��<�k����ҫE�>��������g���O���C�����%͗`f�y��¤�2ˁh�N��c�J���)��+&I��u�T(쌼->+%�u�v�������yv�0�Yj�Vx��	VM��a#���VD�x�o^����Mؼق7�g%�����K~tg2i�A0N�o��Z�<2�%���4d[����#|����j�/J"�D����c�]ж@<;��3ɟ�?��N�bQ�P�@�C�Ԛ�%��T�����A���o������01�r�hgd:a��VS
D��kRҒ�⢠T��x�*as�]&�MK �|D^C���R��j~,d�����]�C�̳����]�o�M+�ر_�����o>W����ǵ�݄��y�sٴ���� �o��-��?�}��������^: ���b�n�Er;ˊ�S�EKY03v-��6tny�.�]
@���O=��}
N9���4�_~��xH*A��1f����ؚe��xS��Rx:z����D$�s�8o8��B���V˅�+˨6*h�<5N5;S��z�>�n��E�|rN�������sR0�ZS�m}}����JGM㹽�Ш�1}xO�~�П�;.��{����������&�'?��p��;���ŕWݨ��Q'o����}2��#��3�:�<����C�����>�k�n�j��W��� C_��������i�T�-��(��8&/i����To&��fB`�Y�X�\�*�l���E��p�&����v�~��O=��s��h���઩��9h�j�A��_97XV�٪��X�M��������h3�U�2 �Y����j��|�B9'Y8��O�z|O��]O���saUCFt`5�/�o�*
0Ƥ�`�V39%�n'v������m�M�ݑ� W¾)����X�P��3����Mt�4b�H�I�>��I�$�% ܭ(�ը6ЮU�70`�`�����dK�b���bs h�	�#僁�a����q�v,�*825�C��b�XA�;߃e�y������3�j������������7�{�/��x%ӡI��
n"V�Le3�J�[�C��fh<���iⲊ�?����&�=���4��4��-���🈰���(�-9a ����U���lϭTd&��P{U�R�1��F��B|xP��k1��*�:	0�Fȁo� �!:�&Y���7�Z�*��߮jdFLA�c���2�ι�� e�����_O�n�>+ry��3@��y��01m�B���k���
 �-�2h��3���o4�����
�j�N�<�u8	�>#�u�u�jl��k~��~����(���!��vx?A�\E#$3|��\ŏU	��`�fXxK��|U�    IDATi��;�����ý6�U��y����K��!�G�Z������{I����I�M�@vh&?W\��u�(���'����CG0��`]���ض˳����9f^PR��7�3��4ߛk�������}�Iځ��}H/q�����b]KB��z��2�tp~���xB+8�s�.W���������g�g��#�dI{]��d���{W�C݌R����|?*,�z�:�����bX��T����G0�Ob�ݷb��Gp����༳�m�����7E/�\��bS#�C�3�ߏ�����TT���Ȃ9}4"$y�	΋/Ə����q�xe���9�M�~e3�_^�����r�U�!ZJ��Q��\*z����R��"�}��E�P�j	�Oڎ�~���߾�v�2�!�Y��p��P^L�!�	�B�O�ga�Xo�<�V�4�N���{��uH] "&&�n�/C�	<��!|�?�Oo���Z'��_���E��"��B/��
�J\P����8���ڵkp��;�LM�����(�����֝�w���ǰ{�c�<6�N'"*�6I��]�궗��:���\ ��X7��l�o8��s2f������Qk��	` ����/}��nۄ���J�KK��<���9)=mZ�g�<��t
6�]��d˅9�t��7�#.���9��{��5`�S��ڞ��T�礮����R�*�Hln��#��p`�AL�G>;��t	�?��/`��6��?��^�>�t�|�~E�?�����N�<���j�{�0���Ѿ�oś.z����*<������o�ş��]���~�����o��o^��yi�����Z4�1]q������ԄP��k������8�Gn�j�;4GAv0O	e���eX�¶��Kr$_'�Uhy6���ҟ a�]u�jO�"d���
-p�W��00�,�����xhK�B�V�d����j����9��[��7����W4�l�\~������werS���>V�m�����c��+bT��É�b���F����*&T��R>���ˊ�g�>d��ޕ�����Ԟ�S���hbt�l�q<6mފd6���yLN�"'�º?|ͯW��3�̃�-g�Y0�c�)P'�(�{tI����M�\�md< 5ށၙP�T:�"a�V�E~+��ys瞈��5�<`�qu��ϻ��IbY�j m�:c9b��$g�����k�[R`��π+�b�	=+,�:gP����fn�
�R$2 ��*�N��IԂ+o�SJ��LS�a2d�&��a F��|�?O^�'�
&�ɠ�l�*��=z�Wi�z�O���:P ���q�`0"}�2�G�;,ύ�<q��Qߞ����`��a|�*լ`�=�o߮g�
�%������p�P	�Ǉ��H�k=�5�x���0G��4�K	]���0�k�jp:&��������W5?H�x�WO-�3.��e�~vp��G1��S�ˀ��Ov&�E�t5�t�#�ϋ��v8a��4B:����ʺ/�iQl�k�>#��`Pίo�.%=!�{>����EAcx+�=j,�q�� x�O}v��}��9V\J@{�S<���'D4��H*_SRG!$Y�N�Ln��&^7��`b��4���g� ��[�1� �8�f\�l?<ѳ�ƀ>�ʩI��*O
q�Ӣ5�@��s���Iӭ�1ڗ�i'n�h�����^�UA~bTE#�G�f���R�A�֙��1i;�3�ћ������̼������Ǆ�	Α�<�̋8xtF>��U�ܒ��u�����
n�8�.y(�	B,Az�kO՚��	=��o�9����#���<��{�$��Zc�x�e�ୗ\����)�Cc��,]O4b�UQ����fj�Ȥ�:����^��f2�^�q�F��Kt)�A�A?����7;��z7��S����v�,���7��_�K\r��9`]��b��l�6��$o96��\,(8��]�54:��{����<��{��2���+!�Pb���L+>ȏDP�2ڕE���X�e-�ص��s
r�iT��;�"
�E$9��.�2ff'�~�Z�8����a�R���ff�035�v���Tg��'w<6ML��9�:�ޛ48��Q��&D��k��q��YVrًٌ���&ʸKA?�@�RǞ^ƞ�/azz�J�Xù��2��!��	��7ކ?��a癧≗��?��?bl�Z|�C��M��{Ʒ��}<��~�clٶ�x�;�Ƌ�]��p�MWa����>��~�S�~�ͯ6�׿���﮽�o��M�8\���@;݇H�n���a0�Z�!!`&�w�}�T 
��V�cIj2�@4�̈́A�O���i�!�`B�(rV i�&�x����QI���FuZu���*��V��66�TVAw�L�����iMX�*����7b|��j�L_\	G�d��^a�d�P��TL�x��˃���w�(��a��y]F.cc7���*��*=X�c�yR6��L"iUp:FJ�;�<��}T!�P�8u�41�
����B�9��I��Z�"�����e��8���������y��{��0�z���kC��/#���P�@N! 4�aB�`����-n�RU�tQ+T0�G��9��?�/g���UVTH�}�~����!yqZ�kg@���d �����DB���A��B��CH��\o{�ǲ�'<x*$��ҝN�X����&G	]�x�m��JeE:2��ł
^<�	�Q�֎���ÒA^��-vt�%^?��C�&[��ڹ>y���u��y|�~{������y��^Q-�_��Y>ļS �\܂GB8���~rέ[�^AmqyY��j#����tH�@��㶙�k���@1�&��P�lvo<`�V�PE��#�d��л���^N��z����x�����@���U�=XQ�r�m)��Q�T���ڊ�q3��$��I��Y��:��ך5Q����@�m�&b��8ӿ����1�Lk��q�y��R7>9?���Q73r�-&z�PSj3�KH���Up�DL���d)��>�|=�ǋZ�ˋ�4I��҉g�߯���qN����4�$��*8�!9�"_�{���?v�ǆw=}W��N���}?K�=��w0����"ŤnTFW�b[&F�מ�H��[��
�/=��?� �g��~��E8��5x���:�|�����q�ӳ8v�(ftJ��i�.ǖIEJŤZ�ҵ���*����r�oøIgT��{6��[�����ƙ{��͛%�̿�y�]z5v�yV2Qer���:
q��i��qg���#y�"-pkO����?�j,�\n�W�n{�nT�:yQ�s^&��*���^g�0Rö�	<��~<��e������I'm���)\z��������j -($��F&�,ͮ�91h���	,;��"��~\s�u���s��,	�N#K	�KIXk�P�:*Ouq�2�)�Y;��'n����!?҇�3�P(/ �d;�F����#r�����w`d|Lh���2�gg��g�M�����l�׭�x���X�f�dM�k�I3!���<-%��5���n����?�j�ff�H���9<��s86I�^���8�<��,N.�5g���]�~��͗`~y��z-n���~����?��lކ_��>��7���ۏx"�|�ø�7���Ǳg�4n�����޻��t|����_����'I�������8Zj�_��t?"� �0�������7���̫cx^����#8c��S��5_��b��z-��5�֒e��-�B
_�*�R�-HIF�lYB�Ā�Zɂ0�>;X��[�ePS{1���ۤ�-�6�E��;�I������A��`�[�"�Jf�&�%<��c���lF
'��zx ��o�2�UZ?�V��������F)I�Q+��fS��L���DĂ{�Vu��2����t-�� �ɓK�*��}t���Nj;��2n�U��5�Q,.�����8��T�؄!���1a;+���{ld����pK
����o�nV|:j��I�xB%�!����K�$వ�� W�z���-�-OΣ5#���l������a�R�����3������a0���2����dPE��$w�W(��B����<���(�h�����സ\T57�?�����p�feM�c�a<����	�C�����t�*�w�L������@�{����Uqޏ'l� qȑ��df)9G��H/��a���n��t$#��j���ǒs^z�����4��y֒rw�V����)Qv�a[Y���^Ʉ��*&Gf�F9P;��m۪�"���Y���Zf�C�&j�3@OƤG�&1�	��������&~�
���l��7!۷nS�{>v옞9�����cG�0�g˪��,y�^̹ R���7Y{��^/�{$-o�՝3��imH9%����'XS3(�2�M����a�Ν�2>��ӽq�VCz �kg��ƔX�&s��hm8�z�%B|>����(��NH4a2��y��>ǅc�E%n����sA
<�+� ��_C����1�+٢�ձؑI�iu0�g����g�k��[+.�
Nپo�[�0;�����Bcv
q�����4�����C
B��0��|,I�!!N<Jߟ�Y�+D���Xs��Dȁ"�N��ύ&ɹK)9��B��8aM�B7@WA�B�I�!j{~��f�l[�n���K(���May9�q�Z�F�Z^qNhT��&�IS��p$[��MI-����^��w��<+��l��ܓU�{��U�Y
�Y�{t�-�
�-K���B�֭݌Z���r�D&�u,��Ν[��8.}�&fg�P*�E�N�鳑�>F�$"%�G�џKh�]*07��X4����ಙ���=��sE�ݻ�S���;�Ʊ�G��!����%�)�b���1V�)�̵���1�r��Z3@�2*�"*�"�F���%���09uXR�#�ؼ}3F֌"���7�����4�utjd�ql[��m݂��<���2��zC��PT�N����Q�sO���ۏg��VS,C�C�Caf�����/ř;�ć>�����H�������>��� .~���|[�l��n���������p��.�G��8��M(7��~��r�ya/����w������7ڦ��^U��o���Ӿ}�m�8Zj���(�Cch������(op׊F����[F��D,x]	C���GV��T5<�4k1w06dy�3���@~�s���W���zτ�P��Th�"gW.��`�
\�X�%�
!�D����W2݉ӯë���LQ���5�|�i��A��c5Ք�k��?1�j��I�WV�o0���F8��*�g��<�Hr,���YоRZ�a>2A�gĄ�*y����ղqrC,1r�됸�-�p��"F�ҁ���L�I��[�2�{��+�.�P�聲�8�=FM>L�N�|2Ą���TmiW�RE�?��A�}b#9B�N]!:i'[��9o��;��pg2�1�+���r��ʄ�EU� ���V~�He��Ԫ���4�d �˩OWRVP�Ҧ����z$���:5|~�|��k��Y`044�f�Dɞ�%d$5�!'�8�aʪ��( �$���d9�#�=�P���dr��+��|1ErW���!�Á4V����Wt9�ه���_���ϖ�Ʉ��4���(�c"J�\	���p�YE�Z"��ő��ίf��Bq��z%F��(�
�~V�W�(����ú��@�h��2XY�2���V�`k�Ǘ�(}r�X0���'$�2����#���f��׼#F9$P��K�cغy�?4����%�#��$�y������M���θ9�XնĨ)i?�CV�Y�z)
q�\�.���-U���J���C�={��Q��I*�֬�nk���#��k`hP��~� �z�|�<��k�Q9Δt��s?�:cLhB�c�� O���"1�&`���HH"c�$�;Ns�/uH$��6:Lt�g`�U���Y����� eF3�<��l�39�b$���^���:��?���t`?y�=�#ƹFY\���:��&�'�tӖ\*YUp�U���֩�t�6dU~�KM�������E9�-�T�C�d|�<��ha�o[�ƹ`��ǎ�)av�7����3������ӺW��{�+d	W��@�}P:,.��E�޳X9X����1�9�BW[W݋t��^��/U!�{��3!t6�e׎2���tSga�<��w���|�S���s15uO=��x�t#	���\-P,��o|-�v�E�"�<��7j�r}C(Uj8c�����]R���Z��+��cS�޿� ��t��0A$�>.���*���<b��iq���F�e�f�y�N��bvq
����3��M �R/��8;��ĺ	�ݸcc���F�'(-�(UP�PD�K��I�1��c��uR%"l�
�ƣp����[й���q�r.LNOi��+�F���їD������?��v?�3v����x�oD���=�~p�5ؽ�	틯����O�)֯Ǎ�_�o�:_��O>��.x��7�<�,�|��~�	L-̡/}�/�x�'?����Io��ʿ�����߹��������E�m#�?H �f�~=�L-n�Q�:4�an�7m�ʔ99,�P��R��2z����+u�R���"#,ː(@n��`�7X�-ᢖ�%M�Ӎ􂙫�Oą�	2�v������C(��h�~�t6L��_�M�C�_L:)�!��x=[��`��N���W�=�v���d`ɱc%�+����a��$Tὅ,7���`=tu��� ��"E�@�6o�S�#A�2��`�=�d���Z�+�%8MH�䨩�G�00U�B˛�A��$�������Omp����޻W�<0ӝ����B�WǜB�`zBƃ��W��mY�ƋgŐ8S�B�u&�b��>Ǆ�V�x<��0���Ȥ��'�7�I"�6�R���&��C��aϪ�А�:r�jys��Zx�J�C�*���&� �``��C/�K��H��wa����#�����ս�ˣ�񼲓d8c��*a�p����[�:ܜԥ�B]���s8ׅ�!�f��׆w8��KX���{L�>�c�b�%Z[t 'V5$e���9jC�^�r��z�>���wW:���S��p0��U���'��9l��9���x%�:ԍ�b�7R�����޺Uά����~x�Z��I݇�uV4����w~p>;>C��S���J�/�l������2]325�������C�|%�a�c�%u�R�'kM+ y�ǯM�s�6F���N�� erأ��|O&�jE�CCBy��ٽ4x�U�C��w��ã�DI�d(�0x旺b���s�[��U��eA��\�׭Q �s\�@&��gıd���I� �>�D�(�	��u�*՞�?odd#�>lߴ�Nzq��w�w�C�:*��rD�nz�x��{�R,#lne��D�S���0��ƹ�<&���a�|�&�M(J���f��.�T���5ó������A^��T
��:;O;UPJ&����GaiiE�4jғbd��g� A��_A�+D�q8���X t�yM�Xx���ÅK,~�X���7	��BR��a��~,�&��S](J�_�h���y�F|�o��w*^~y~p�����S��_��!j��J��V��?������%���?n��O�ҾC(U;��_�q;����_�m[�┓OĶ-:Jx�Q
��o�5�^��/��1�H��MU�X��e�=���C�;wM���y��ݰ�}:��Hf��g9-�E4[5T�%A��0�q=�mX�5��KR:='j�%T���بI�~p o�Q!�X�����B�Ji�l�V��X*�8L�1dq�d?r�aD:)L�Ğ��bar�7��w��y������g��O�w�s?"�<�sv��/|�Ӓ������_܍��?o���Q=��˸e���    IDAT�gw��}���l`��@��������O����`��?^UB�g���S�����Mף�cp,�B�{-d��!���ΘJ��>��Z�$Ӧ��Y4��U_�Q�W$ض� ���η�2��7�Ʉ���	�\|ʕA�^���qm�.�hv��3�J�yJe(BHE�-�7,�*�<�	�D�W<�RO�-ͭ,�`[�]�d+y
_~����}����NXUiS&%��j�OAK�9%�`i���4Ң�M;n~�;��@�)#����CA�_�ê��vYu�S*K����~�<��(���e2ƍ�;6��w��;Yyu� 8AH<D\	�]��?�d�V�O��Ǫ9��rf�;
|nL 8^�m�T�'�3`1<n�{v�\��&V2�f��TV�?VA��4F��E�+J�>6�*�x��)�n�dp���-8�Ӊ�#1��!I.����"�,�)�$�$n�1���BC��Xg�s7p	�K�*l�V鷷:ґ_����ܞ^x�{��L�e�a������E����������P�1�,��w���0A��\�<$MҨ���hx4������a��&�UYÞ�]8�C�]�N�(9�?�Jhpo��}��;�TVY�P#(�9(6܇>�:,�1��f�%��	#ׄ�ޥ����.��;���ͫV����=�1�
\��{L8^�㰺5�����ӡڈ���H�@k�$iI���~O�ezct&\��<�m۶mul۶m�NǶ�tlw�a��}�of�ܙ{~W�U�N�]�jX��?l\]�BTƶe��M'����KGF���#��Z�}
*� f�Ks����o�Ms�?�b��%���iΒw\���@�w�)S�����'V9�-�V2�h{\�B5}�����&a�.���Wd?�u�Z��y�/w��n�{(��X��X�(�g�n%	F?��#�H��������GQ[]�[�js�C��� ,�%By��3šp�Y�Q�|���B����qN�^ɳr�<X�����W������2�7i�����`LR�1u�y,����x����s�#<��������P�N�aXA0�Rf�����E�yjy��ۨ��Oz,��=ǣ��.j�Ұ��墵�r5�H���z�b�;D�޶�c�Gy�Q:��	��$������y�4U���q�z���,��d�.��b��\�����A�t�>ܲ'f���sө�8��iR�a,����:Y^��Gw���^�������M��j���k�mWz���޽�<؉�`�+K?� 0��u˃���w9.�ya�`/=Z����|<���F���.�b9�a��U��o��-ɩ�63Z��ۢ���
8�:1]Z*�ӡ��Yf^CH���7�#W�?���Q��a��a;����|0x���������i��U�Hپ�m9�e)~S��:���)S��pI%e��	ul�V�qs���sן3W�Tr���#��,�]�]������W�����
%���>M���^Qлe�W������)����W�xv��[���/(��ɇ%N\�ւ};��MGBS0A�)�a<�؂z��ʳΌ���E^�"�P�n���t�!TS��DV�|H���Ï�ͺ̓�h����]�yX��?afj/�JM2�$v95Ra��UG���d�F��v�ۆP�F����"����e��t�73���-|VL�gS�[��-��Gk>��N��$���W1Ibv��.������r�Q��>4D5���|Q��j�h:\b� ?ݼj���i�J�� ~0���3aB��n5�j'<O~8Pm;Y��ĥ��yO=�eP�_���80c"��XQs�]7����f�tEE*�����=��E,%����\,3 �9�K�q���#��&�����i�ˣ�)�D�_$㋵�����3e�#�Ƞu�@���S&���#4��.�n3�X���X�v�(�Ii��k\�MZ��'c�*���[TV�6>��ԇ��N���P[AA�
�~�\��WV��|yDf�dZ���Qi�aE..� ������߇i�}̿������X���y���-�6��a���Ggq�.�~U"�Ës[������X�������i|���_�4T��O�r	gPB���i;���"g�Y�ff�¶i����ؤ��w��{q����r��	u��g`��""F����^s��Jz�X�`�i�+Q'!$�x#�I�M��*,�nH���UYn��0��V߮�wY,/��^�L �!�mvKª]lJ�Y�m��E$�,ٯ[�`G�Ds�L��������"�_�J �ûA�nL?�X����P]~������b�G����L����K��AU��f��D�HV(�a�ǹ�]{�a.d�Y�"+�O��;�<3�,u���Z.�rX�ٟ�m$3u� �]K�A�{}���f�Z:tsV'��Ƅh/Ѻ:�T�E�Vꇗ�-s������վ�����*c�^P�|�O?��Z8�3Y	�����݀f\��!g[�l���5����͋���O��b鼱�\(���v���r�W�X��I/w���q�������]�ȣ�Q��f�&���|Bo�{��Myb�R����������`?�2w%Z+��X��&=�l��5}⸝.��ْ�4�Ua�V�*�=/��wQ���q�OG�:���&[Y��:�*�{%�'+ŉ�����p�;�Ĕ-N7Z,'��}h��M±ɮ��.���]����x~��s"D�}ٱ.B!~��D� L���0�jX��}�{�jGK�D���E ܎<���5��=�� ��5�u�ⴚuR�+�?h�A�:w���9
�|Kw��P�W�_ê0d!��#�mӝ�X{�� ������u�m�_,ˁ�If��Pm��=��ӻ��G�����i�z�ƽ�n��Ճ�`�QG��Ͻ3%������Ԍ+�UO�'ߦ�2z��C�u�9�"'$�ՕB�f�$J�"�6-�uƝuѪ�4�k��4�ž׆�b�]���~%I�6ߚ=g�+ʔ9�eA��:�v�J3�i��}k?���*4��hL%ʞ����g&����ѓ��|qҒ#�M;.��ҳb'΃w��RSFҤђYq̤�>�L��f�ҽeɪ�8I�b�-gƝ�Dщm��CyA�e
/�B��f򭝡5j� ɞ�� 7J��R�g�q'�L��~�Ъ}+I���,��]���,zR�y#�!'a�4�3�U�~tO8F���ogc��/�<;�	��f���Z">�b���<��Rd�� MYy�a�8~�9,�1J4*k����d27��F�a���ds�+眚L��C�b� X,����f&T�l��2��9;�_&���[Oy�thPP)䛾��>�뜚�c}	��V6a�賂"S��V���lث�"�af�h1BE�Ɗg�{���9�x$.:��/A����*�����|[��zϒ�^D:N�(r;*��<F,��r<!���Ţ�@(w�e�5U��=L��P��.���}r�yƧ�����8E�<�g{�X0�Y��V�=��6����2G�"ؘchà	�R��ȩ!V����gn}|�{�?a��$���'K���hL��n0�1��K���}�?�ݪ����%�$�bw9�F~���)d(BFA�CzT�o@��;�!�=9��7L���:'�2��`��'�>�fo;<BV�b��� ͜�g|E|2dY��GA��B��P.��ui�����e��t��EuZ���Q{Y��E8���e����D�����1,3P�V	���b��q+��;�eA{�����^�bH�!�y1�;�@����3=C�K�}Ō��Cd%�'xQ��k����d_w=*�i���QMHH���Jb=�x�dB�2����̑��@*�v=RgX<PC�H��S�wk2a�x�@��YO�x�B�"�-�Մ���M�i6}��r�ïU��Y0}0S�BC�?�*Z,0�>�˝�N&�b�.v���]EB{���'�="��{�sh�s��7�,��x�ґ2��A��r�Ә�A����6��8Y���X�x�w���Ϛ�.So���#�vc�	�嶃|�G�g�~	UG{|���5��?^VyoK.����Z�%9�L���{�UY��{#J���|?__�!��)��)	_��^��4�����'C�Z��X�Z���nH.���I5��μ!�:�Ha���T۹���As��j�ӡ��-��P�U�
�qB�C�~�k�禐.��ʃK�j���l���\����~"��!FI��J;�����go��t׽+o?���44��Y���|&��9�]0����?2�����aV�:�y�>p��e5�#ƣ6�Uh6N�?���s�Ѿ��/��p9���Y��k4b������F�o���"��"�%I�RʸH+���p�@W�v�eRlYM���S�<O~������uԜ���$?R��ּ�+���"{����'�/��(O�����2m���G�E�8�����[�ƥz�Ʒb��
�������(r!�*t�
tI���4��/�q�:�R-�1�2�<Jv�٫Z5{�]7k]�0�صg�0/-��m��ZucƗ�ބ��	��tf�yǖ=:�/
�vRc�q��t�� �X�㟹��uڦI��j�2��Vz�l(���X��ڱ�L�W�)/]�)Ǚ�n�=�u�YV�ī]<�V/����,X������r�Č�<z���IO>�n~\�n;�S�i���q��
�D�jԬ�Ք�^�aӉ�쮞�˰;r�F�i�ސ�M:M�ű�Z��8����6��-*�v�I�);�?z�oZ���a㉕0�p��I˩|�?�ѭ7]�]̺F\�휫��4ؒfa�b#6�OB b���BI��BCah��2������
I�QJM���趠	�k&ӗ��wj������i_�ZW�bLb�@���w�<v�������wE�#�0��ln!��i�A��u�$��c�#�ܘ��G.�B�[S��m&������5��hlW�"���r{S$G ҥp'q�W5�Ԏr�����G��b�v�o[�f�k='Ilid���W�	�c.��<���n�7��i g��]h�{�&�7�tQ�:�`�%ލ<F iV����q�T�K�6;�S�n�h�+��h�F<�eT�\�{�M����YR��(o,n$$��m�L��8^���	��]1�Yx���S<[������?����{�}�Zh$�c��G����c�GȎ�UBt�c�2��q[w���t6��zlF��S(L�*B%|�ez�3�#�ӹ!���1�oBֹ��l� q�������j�et�F�I}zl����a8J�d��[va�wau����}H��V�̆<!`�8������y �X��Yq��0m`�'���Fh�'8����/>g]�y���U��cTt��64�M�W �or��\�z#5��O�bN
�q-z'��S��"�A��b��>�c;��`X[������0ץ.]��z�ȥt�(���Ĵ�+�[oc���$�>$���c�pV'6����pk�~���T��	aV#�ü�W��i@5aG���_C,� �t,%
�Fi5����o���(������0����N������#���ta���	����[��c>	XFc{��Fܫ�)2'�{�9,��y}hV'����G�3��N�Ukp�����!p㡽6��钳���\�򾕭/���여�M{����{0�X |��c`�|�<۬"ɝ�_{C�����V�^z����?/K�懨�Rw(_>��!"���o �ˊ;|'�Ͽ�~O��������.��KV��rCNB���>�1A��P�ȴ�g&6mMeâ�!��<L�����b���8H���ǂY��EU.t���K���+�ct��A�/��F��S�]�,�4����z��6g;$��`ɽI����/ue��=�q���C��V����9�Wȿ��8]p( ����z6����=��}�v���0Y-(G����X�/T~�u�����s���T�%?����<
�t����~߿o�����<{Tص�P$|:�yB����Z;),1-���X;t������ qJ&Y1�YuW��ڤt�2,]]B۬��uMG�!��]��e�-��j^C!���Wt�o�3ow�R���ʺ��ͤ?���Q�[�
;��`��]Xթ-s�b>��f�)��Qv�'���ӝ�lt��K��լ�Q?�����Qh���}���i�ֹ�3s�꫟9f&�աks����ͤ(��g�ʼ�TE�y��jh��N28ȆF��?P����eW�"��&_�����:R!��{���G�[��P����ﶍ�,C�6��?�>tN���!9ą�'�Ǽ	G��Y��w_��g��n䟃w䩺�$�#�+H��G��zͭ�
�.^X���n���{�En�Y���n ��/�=���u4\K
��]��Z;6���<��ֆ�ÕP7�t�/��͍�	4��gH�Cf��%�M(��n�f�S<"h�|��f�� y��6�T�U��j���	��s{��p[H���c�?�JD�Cݫ�P{�J�%1���X�a:]m��ÈK�id���=�6�& v�����L0�%������fq�x��&BC��{���_A��ұ@��V�� ��`�bЈY��(��׌$(��ER�F���-"��@�)D��[[٣�̏�Y�e��~E��:�Tx����U�Jr���}/j��������%�,a�Egz�̿!8�����s�lݦ�?k�1wN�y�t��Ï�F�I��G,RQx�}
`\K{
�.@@�� ya���!P>!np��P���m���?ɦW���N���Ģ;�=D?x�l�B�L�-P��Զ+!�����{�@����B
#���<$tx��v��`�z+��خ�n�����!J�#ô�|$�ZA�aГ��S�c���O���y���q3����ʠ���샰)��B��t�E����A�~��#l��_����;>��:�v��n���h�-�� c�xi�Q������Y�{l��S���b���v��=��/'G���s"����]���i�Tuz�, �fQPX/x�6���RK�٘���(	��-}�r��1��^�9T��F�o���>���}���B������uB
i7�}� ;������`�H-�L&1!��]���dJ��0d�3���(��dc���O?	�؄hP��1��Xw9��Nr�Q�8��b%iae��-4�O�꽁z�4���y�͢��g)���w/K�p�K&���ŉ=t���yE���]����k}\�d��F>9��\���������}��-Q`O�9l�&��_����?�uk� �0��?��l��L�>��F��tI���S+�+�EY����s��P�X�6W7�\*������;�.|9�t�3+�sNX�����nS
ٻ�뜳V�U�5�=<���(:sq���ԩ��ڀ�|�� ȕ?:[tU�to�Dd�s�L�M�Y4�vo�I��>J�J-%)��A�b]��o�ks�ᦘ���K���{����[����AfkiP��.j�AP�=��a���v!�oMtU2a����K�'H��97����p�f�׃�_��O0���s~X>` �����%��
����8i���\����C��.c�<^8C5����0z�>5%%š�3�JY��Y���p�mE3z�:��C����Ii	�c�ʦ��Iמr�R�����7�;���oA@}����8 ̈-��g��6֒q%%�)��A�\bf��塠�iǆg��×�B�k8��u�[�q�ž��樓����,
~�&�ʮx�07+h��rSQ�)��@���zD������P}�I�>G��2����V&�)������t��|���ث#�T�t�
T��܇+����d˪�LH%pz���{��h��4��Р��k�r;* ̾\`*�T����.�6\>:ȉ	0���=�f9Ԉ5���^��K1L� ��
.ڤ��� 2f��/�堜��b�a�弖Dj�q}�4ّ��;T ���68CP�+H@��8'�e�K��E姠������'��K�7��l/�Qȃ�p��G_�����UϪ�D���R�9�j���u����ԙJ7��� 6z��T TH^��~G�	޺;�N��vv�j6���X���[���@�bcT| kgi�� �iy(<e���4�2�;�(]�a+Z�>�4l�����vd���j+�����;>��n�T2>�z�̪��wY��Ϸ�*�/r�]fPX"�q�( d��Y��J���k+so���w���6OOX	�z]�'ྲྀ�0#��<�J8�<$,:xU4�r���( ����e�F�ܬ�䈇z�l?Mx�|�Tܑ��6��^�Y�yL���-�cA��8T�	�}��K'�u#�w��ܱ;��a�u���ߺC��i�zYc���+�}�G�F.A_��l�G��@�/� �H|�L2ar�3�ƭ�o���b�,���ʬ]LQ�-f�߯�'x�����|�'���;��i��<IU*��Uק����g��FJm�#\DT}���%Y�'e�����3�/F�i�c<;��7����ݎ?�_�~��o6�P��o_'� �9��=*-�ħ#�~��y�2Z�'��.��Q>Sr�,��m�1�zܺIu�,�Y?�jR�)��o_�����/��."}���P��-��k�a?p�=��rol�
��Y�iN�f�v/*�D���.�әY��7O�Q��s�K�Zsi��n�y�SS�ҩ4u�Y��f���=o����uk��a�Y��(K�l�"h0Ð�"�x��h��&S'��Xle]ӭ&X0V�M�O:`���\W�D�轖��.�pA�h�xN̨m�~�J�� U�g]��6��|ŋ�+S�|G�"A�����S]��N���\]�}-��K��ɫ��>�N����Oj*�����`���m�1Qm����8���h�	�,��I��AZ��B	�K]�Y(1����`�BdkSڞ{W�|� �A�.�YLq��yF�g� ���� �PI��fl��R�n8�+�?o�&�����e!��1lC���w���*��i�pD0eԮҍ�����:�:�A���U�ӗ	L?�\.�'�3$�o&�#
cSj�Ĉ��@.Kt"��P�n�4�͊=�W2�?�ZѩÑ>!��}P)SB���T0���X8SL`�%3*�Z!�)��r�57-����p?%@Y\5C�m<n@�1g��a�a�u�-	������8��`#����F�)��x�bCi���Z2�����w��*�l7_rΤ��0;[�KRO+p��y���c�9�6�$�����ЁL �Z'�	�S�;����q,� گ/��a(l[b@me��Ψ�Z2Vf+E5'´D Y�1Z�E�-7AqC�y�|��b[�a�1h��r���H^$�|H���
־��Ê� 12}�22d�����N����{�F_~<�D����֠�6OO��\��1��c_Qi&�5v�X���O������R��'7���|��8a���yJh���,H�Þy�	��O���%�3�j�a6��SwGg)�<�$��8-���j���a��:���Z�QL��%Z�K =��ɀ�'<�#\��0h�!���j9����?TMbq;����6^�lQ�/!^�9�DB������e��ҁ_>A�=��-I��?�W��N�nG;����ދև����"�y�[����G����w�����Y�oS>Wes�7f<�GV<��c&�.�D�Q�������C>M.i�5�|�f<��N�"��s G�w&W�̘�Ǌ�DN:mZ˩��$�ŭ��e��Y�����14�7�!�g�������d��t+�U����q'jZ'�������t+	1��G�'U�#V�u��Q�z��)8QReի���ž�TC�c�u,���e��J���^�(�,j���\(�U�*Kx��h���8o��f�-��e�ַ��b�Q�H�,�J9�F��|(���:Z~��Jv˭Ӄ�t�2ɪ�l�Y���ۢ$@�̈�eu����Y���0n%/�{���֮A�����j�?u([����:¡1��iX�[�9"»m�d[|�f""�'kW�>-���M�	E��x�Sԝ����6�)���/��=|�5�t�F(��1�}�A���G��8P�������b4�P��x�� @16eX��^�Ÿ��aA�52��njfԣ����f��Kp��1��
��ǀ5��e�B�|�׌p �K G�XL`�l�.�8��Mc�}G׮7��~�\�Aj������M��BGM����e�$K8�~���r';=C���b��u=╇Y�	g�ŊD1�����Mq_�y8|ȩT Ao��]�����9�D �f�T��*47��J���(:��+`��B�-��oD ���(���$H�/��U0���X&i�g�[r��1���!F�2B�d��6v�հs�?!y�7E�aQo׸<Z�c5p�{�{ֺ֟��|����}3����+����B)�~x/���j=��#�l�2A�m�G��ξ$���-��#�]�UH�V%A�qz�O ��(�M(���a:���J�#��W�x���Ё����n����G��Ү�h xC��u���O7s�?Sߊϸ��	�������W@ҡ�����J�lӦ������P�+��a�~�v����������hs�;^�Rq���/PA�?>��e���ɮ}����c<I��������_�/P��x=����lEd��r;��.� �GTy�j㪯ɥ;.&@SQ+��1�b�t	B0�Y����f/k0���P���ݾ5�����^�ư��;�ֽo��wf�8�diÞ�& ���ҾҼQ�P���I����ǰ1����tN�}Ϟ\��V�k�L�8�8��ުEl�R�c��f9CoF��GX�>�.ĝF9kg[�[Y�(�Mvt�v��#�@�8�j�c�pQ�������:�*mip�s�o�M��¼F\����t�6�P�,XCM��N m��6С�y�t%rh���<�6+�^a5�R6��~pF��"6z�y>;��=ـ���:�ǽU�ɮ'�Q�(J�Y�v�8$͗) w=�m{�Kp���v�O��B!4��_�/��"[;Ǐ�	�z��|�9�a"��o���:���q����\r;
����$�pS=�T�dˑ�ʸׯ7����Tb0)��`	�'I����β���'J���c�N�@��9�{!@�X5�v�[�e�1��|$�%�Bc�1 iO�R`�%�.�!T4������R5r���v݄�fi�@�w%�1�t�Γ�Y��P��Ek��$b�߶��S#��sX�+�'�l�<��~�;T�����-ũ��*	�]8C�����:�#�\�W4��e���L��̱���PM��"���}y(\�0�g�<�)x�;/"<�ꖮ�_c����ς8�L����?C��8b��Tz�G��%���~�{IG �ņ�[p�-�3,T(����eY(,#��7g�r�ݲ�p����V��H�����b˄O�����=�i��t�V��0����|B�mv���w?PUcYf�^B�}�W)��{���[w_&=�<���5?Ze�����3Os��;̡�ӽ�kOH���{
����X&}�%s��g��vc�NtӄX�謭]o�o�t�ܑe�����IF���ۦ�s�D���oI\���AV�%�	��O*�WO�1��s�i`�|9�;�V�{=�Z��(h)ע�Nc��Lt.�Y���6C�o"c�5K�Pj�L.:�<�I3�k� ��Ѥt0�R��lF
�n<9��ƣ^!t�W`8w�2̦T�|�/׊�9
�Mʁ>"<�R.W
��[;�,�4� �@x���V����[&(H�7��DOJ��{�3 0X'�O��e��!�M!�Y�,��S���Yp�E ��\��&�M� �	2 ��AR�T�U@�2j�Պ��^ȢZ��(J�����O�vk�2�{#�-�ta� F�a�/Q�p���.Ƥ�ñ���Rh��/͈)�Y�j~k/>�J���K�RE�&(�\�dy2�f!�ؑ7�T�ڀr�0�˶	�V�����#���s�?I=���C4% ���u�B�J��}b���!!�2 �9:��3v��� �dix,w��޼�7'��o	�t��*�r~_db��
�N�(��wǌ�#6=�=�N�A�}�0�1!��]�GR2�P��覭�#��{/�O9�$��Q^���\G����� ��g�܁�	,O���ܭ��U����q�b�-=�7��y`	�"$��&kBi�����R"(F�u��O���?|&�q�Ʌ���t���=���s�R�O��Y.I���wT?�u{�U�����gg�®�?7�o0�ټ|� �+�u��9���n�]�l8�%[[�����l�S9z�5I����[1rЌ�.�������n+^��kGvk��:� ���`�^��m�$٢��fK���&��dev�)m�L���9�4�j��ra�pL�t� 쥺˙rH�C�<Ny~m���7)e,*���M�,bm��J�X���.+��[e�nW2����g}�v�ܠ#1w�jYM��b�f	7$Z��l 7�\��S�'-S�D4z�r�(~-�V�2{�Ie-:/odu��ٓ�β�*��,^���i/��	.E��K<Rk��t���Cw},�S����P
����b9����^�#�^}��&[,����G�H
�
 3�Ϗ�&���Vt�i����=�ӕ��Yq���;]�\.B���҂L�#	f�4Q�/>��,�Z�р ȫ���-='q��^9!�P"@l���NI��)�=j�4��2�.& �]8k�bfk�/1�ѳz�gˉ�N ���B�Jk7ˍ���ac��i�J%דd��h)���bt��H����V�jA*He��.�1Ĭ��}C��-l ��\�����H$!W`ݯ5�xa�;�@I!�Z���A�Ym��]�7����5�E�y4D^�豕����l�ooX=����Iť�C{���6|6��'���篋��2����Y��[s���FA��b����s8'����w��)�����=UBG`?e��Řq�?� ���rl[d�mG^ Kh�2�4_m�N�{��I�����^���ꫫȺ4�-��SGJ>2Um8+��t���Wq���=�B�=��+®L�cU���br�.��yL�е�6� /!��:S	6,�[@7�y'��,��V㫪h�`f����<���-""b2H�����z�z̫��I��$s�0���W7�H#JW�����W���l�")�R�W����C�m���M���9y��)+��rᤃ�
���rE�3F^M�
�U�h�r���@laa�9B��Mnؖ��a���2��a�(�4�m����K3��{� d�e�#�X2�j!컇���)�~U���@�ɟ�<�@��䐵$т��Qj� sd��H�ͣ��Q'��s�d^���� �i�U��9��4�(��?!� �Pe&b]�X<?�ㄑ��@~ɜ�
��uX8�����t&b���(�D���'$�!�]|J����|�,�A�YJ�kǈe;��-�(|"t�M`�`S�*��&d�ٖ�&�}�9�^�l�TG��\�@mM�a�I�:��2ؿ��7����5�a@B�qO��X�J��1��qFވ���X�|�УE�?|--O�pEc�+N���ߓv�Eqm2
^h��v�+
�J�-��r��z�>�$�~Jϱ��-I�j�������Z�|���'��x���(�2�Wq��l��Ϝo��E�U��IP����N����z��e&�:���s Rue����l���H�;�r-�5����N:�==֠���%9󥮠!���0�7xJ��q�e􅶨��ڠ�����!�ꦟ�n�Y7/J�PQ�nm��=/JS��\��w�+��F�,�g9��T��ӭ�E�	�9t�(�>�9�-��L�&G�^�8<����������}�����TKm�4�m2��ܖ��f�uī��Zl�ԣ�̔�T~�k���XEc�cz�Z�aU�����&�s�}#0
/fi�5���]�[_U����Ɛd���۷N�$l�g@^]㨐�Ț3c��u����!��U9�N�s� qDz�8%��E�WB�y?ȉN���'�=�ɤ,Gi��)n���GL�����i��-�.U�eN�2|��	_����F�u��Eօ�e�!xBj"ZS+\*&��׆[�Nm�NbzT��mh���"��n�o���MG�6A����4duU���!c�������a�g�rS��8�E�g���dy�=�C �IS�Ek�% 0l\^A(�U���7�Ma��<~��dn,<O$@�4& ��\�2���=�>M�%��\^9��7�����"��g�>���'���[x�oӬ�ܟ�[��ϟ�s�e�K'��C���	:�9��v������49��Ei6+��`���/�j��6�#�����|Y�S��nssO�4�/k�m��V�/�պ둮�k��+�r�5<�Ҳ�J_%�)3�l�+��L=����(C3_@�.��d6�Y{��6�hJ-9ԍ>�"������\aq�UWZWݵ���ϥ���Ί�KA��d
3f�1�p���#sFF����f#[�N��f-������y�pR눠MO�;��Z	V�h�M�6�N��ծ[��q�m3;��|�"٢���&e�;g�;��J'Gnp���RH:e�h�����d3��li��j�	�A��1������R}�<v�Ȝ�%^�����a��	nM���$-�,S`��~19Nx���6{ь��:�1'���u��>����#9��l��� �����:ZHb��P��@қD��s����J,��� ��������������:��:�ȟ��	C!�k�%��`�,~��E��ʙAr5��u��cw�^:��8|2�c-P^�\u]�>}p,��`�{<���E��	��tc��s����4���=Et�z��<���_��߼�)n���r�glb28~v���ٵ%��Ő@b��XjC�\�������l���քO.ǜ�*�l��[��\�v�[�>I�� ����/����~h��r���u����I�Wb)Zg�}.uzH^�:�	ǜz�E���e!̟�4����KiK� k��x�E�c�����o}N�/�/u��S8��`���U �2Y����V��_^'6[�E�nj�33�|�++jqT�;y��:d�" 2aX�q#Pc_n��U�5k�<�̔A�"�Ӈ�ϠI\g&��}G"�5�ޟɉ�.K�����>W�x��aV�?�!@�&�'�-ѧ�q!��f�=��W%<6g�X �Ѡq�!�~��T����M�Ɉ�ZLJ�+C��N��5�M��a��{V[����8{��?�� 	K�=�o�^k�^Cҍ �R:�����?�_?5z[�[	�>z�)
OH�9}D�|�w������`
ݿ0��m�]�*�<��"���p��mj�bwο��ZQ���\|����%k���#�M�)K�q�z�춠x7�.K%��"�'�l�ƺ���[��j5DH�	l �V
-�(��3���Ç�����2�YԦ�ӏDo#?F���yd�������!	���ޖ�C�[MO��imY���.p{�<�/=DצV~������rޚw�{
$��%ޚL�H�&�5���a70��TcƉk��;zZmkmkןpf��r�̫m\t�S��q�j
/B����7�ѷ�^c���bL�����%?������rY��e���N�{|A�N�{�n�l%5o?�uk>ks��y��tY�_|a�?ވZ�>�u�R��Ͼ�G;ט��[���a�q��=Y���#�0�]����h���/]qH�D�)v�Vk�g3t������w��c6TѲ0~��P ����`K���ʽL�t_�T���g�#�O�kΚ�(i@�k�sԒ�r��S�~�G�&ayz{�$~}Tc��HU]mn��N��i�܉Z�^,.��M)Yu�bmC2�?��Hh�f��9�Va��NrM�D�lw>�6F��-ʽ{WM�ʀ����1��Ņ�ԞZ(�ڱms\�R������ϞWk�2W-�����,C���l��ܮ�#j���R�r�c�c�	Z���w���l3h����BH�݉q��7��*��H}���ˢ,>=�&��llDM�f��mSm�%6�,���� �!m";=,�N��䲻H���ԕK��=������k��TB���zk�=����{HA��w��P���Ï�͞�w$"V+�c,��\��!������c�q���{o�D�ԓ�_����?����#��ҁ�"�����/�V���n{s���A��:&���ct���������_�Qִ�� �y��
bu"���PK   �cW���/�� Z� /   images/d3087b83-655e-4811-b17d-9d66f7a3b2a5.png��US� ��%�[pw� �5�;��ap� �	n��;���������}����˩���>�j*��(�(   ]^N�  �  �#!�'bh� �T�JI��KIQ��9[�:X �9i�jz�K�ct�B9�nyg`q�,�"	2�Rp����+p9$�)�-��_b)���k=�zCéy��0U�����M>���ô�Æ���;9 �I�Z>�`�^��\i�s`���1 ��Y�"��ҥ�[��#w�U׺�o�11�S� )����G.�+�9R�Z'v��.�@+�R52���x��t4N�X�i�1`{\$����S���4.G��?�b,Wg6������"�c����Y5�G���Ǝ�g�8��1�����̖�?G��kk*�K+��T~M�N�U�7�'�5.�<��>0^d�tx�V�J#��C��}�2��s��I�a}�o~1>sǞV��(~1IUQ������	j���c�����4�|}�t��v��t�X��`�p���r��{A=�%9���A�������k�
;����մ�����gH����*3�9fL�1@D�K9 N�s`)c?�9,�Q�	��l�cU.��!�/�<t	
_��va8�x"qBTֹ�h�3�䮛X]) S�������T�h��oO\�Ŏ��9�H?�d�a�L�&�xu��}dް�Xp�_>G��)��h�o�Mu�c$W�ZB���C`�9P��]�a���]D��f1�C̮��$��B����n)-�>5D�&��#�K쨑� �J��!�F.I��i"�������,�oF�~9B�%����8�C�Yu� Ef��`��-⹠�#9��.ow֑"' b��nյ�cBQ���}[P�D�$�
��h�%�֪u�C[Z��;s��Y�AQ�,��ٴ#�#:�g�Ѹ��B�&�tB~4�X��\�ߜ͙8�������~,�}Y�Fu�+L "���c=�|0a�E@9�v� fo���k�y�T[c�A[���rmd����޵�?��4+!ULA��<�/��EBWaEbE�;��-�L4���/DΔLC�jJ>,�O�[)r�aS�m���k%%$�����UZ�rE�����_���l����1��:+��F6�}�m��|*��h��eB��ͨ��˸�ͷDI�Oۚ�]sZ�MG��_�'J� KMP�ܓ�9�7�7Q藤F��ָ�^���ߘ��Z9�ѕ���j��'��b�1�r{��M�MM�M�B�N
�s�%���*�uY�YE�Mk�������b����He�6�fN�N<}�}C�Y�0��y�xÈi�㉽x��x�x�y�m��Ŗ$���O-�W7+��Z�E{F{ z%��N��.@�7�i�>�
0�ա����ht2��&�l���{A��E4+�,O�9��M��K��s�ڴ�;�������V�N]	�
1:9�'t���u����8kV�J~_S%k�2Bg��wSs�OKū����<3M��d���	��ꑳ���<���Rx��dsu+��O--�zMgY�?��4D�D��֙�+���Yfd�F��o�G��֩ʑS����-���!g(g�������K5�W2m�&�.P��Ѕۙ�/�)����������ƶȑ�~�v��_��i�#�p�s�M�����*��y��Ʌ����f�W.mN��v~d0�Eb�F�����u������k��#�+��iv��j�J��C@����ˆ ����z���'7�2P=0-P��5���-6&>u�	�ktq�_���eFޗ�������eT�TsIK�Wg��6�Y"�"e��anR��b��(/�l ��������H/�Yj���q��8�T��~��`�d���0��$��l ��V>�Y�w�w�Ֆ�m�����:&��cpx7�e���|B�
aY��칺�������'dNdD��+Iޮdi�݄!3�����o۬+Ԅ��Ha����V�3��)�����%?�Т~)�9]�[8Y��-�}����#�"B&����q�+u:H�d�.)���q�X��eAO_��ZEm0p;���0��{���}�� ����v�BQ3=*��Į���X"/:31;�8��~�n����7��6�{(ͱ
Mr2�9&^��&�x��o�4Tm˺�8�~�B��L]Bm����¾*H��Ṿq�����ӗ��o�s���OO!�ê��K^N.�:{P���]�2�o���~?��@7���K,':kb[��Xj�2t�t�H�W������Ӽ��+���_2@���Lk���ĕ���U����8ue#ť�� ���˯����v�vUK��i�u�S��'��'b3�Sy��]h�E��ʃ�b��`����1��4h��׃]l�Y��v}MF��^!���Dyp�q�_z[:$�����������sY�JU.�%»�jre������a�4}��������Y����0;�I����\8htu�<C�ȵ��ө��r.$�q�'w:W��Щiã{u���t���������w��)���Q��w1�K�}+қ�q��X�yCaF�&R*������f���������|����K�'�{
�g�|��4�#��֠@�٠��X�g�����	:ֵ	ߖ�vVvޗ�-����;?r�:[���/����O�O�}�Ke	3���2A��v��wW��D��~��A)H�����? ������ge�pY����W���yX6��<XJ.
��3���.��u:�IF�����^��w]P�CjAg� ū�����2�=u�~�^��?����  �����m|���v���q�?~��������������c\8�@���W��Tfz���I��>f���tn�X�7�sO����훠�e���APn�u��[�sT\3�s��e��s��R����o>x����?��?��?���A-��uz�I-8V�����M��U�*��/!�7/��?�B����Bsڇ*kB��S�����Bwo	�gG���6�R������C0L����/����8?��v����2��fjU�s���b���}YU�������_��3��I��`�0����fnE�,C���M�{Y�<#RSM~�����B�|��O�m�������bu����c;���x���>�[N�V���׃G볯���榰ѳOUsZ�>+���i����zn�4��F���fͮ��U��c�[7����S���y����M���RGQH���d�̱,�Ie�������ᶵ����szm������������%�����������c���A����}O���ŏ�KϚƫ��'����Z�U�p��j�P[c{s��1�y37U
>�G0Q^P�^�?�>X�(�>��V�֕h��*��!�&폹����O��ſ�K�k��tT��|����;��Ck��e<�Ҵu�A�SlF���-�����'�d$/�l���=�Z���ׁ�p�/Ϫ��ju���(jۯ/���έ��0(p� ���@��$!;�P"����^G�#w@I:gV?6!��"���_0rBFKK�`�R�e��h��+����O�p���D6$J���*�Yb�.L�vq���@X9��U��)h(bo��&�7�.���h���o��g'I �����W~�	���p������n�^�ˎ����xȅ�o;�GO��8�k��8�u"B�rC��]�o��t�A^�ܓ���e==�sXD̦�˭�G�q�o��Y`�����(��an�JiBi�~�n���-l�J1Z��'��шp�t;�@��m �R-E~Ҋ@������I]1��{2�Ñg���pB�(ٿa�+u����\�G�������_]�z*j�.ʙ�//����id|,~��X�/9�v*.����G��xױ�tC:��Qj��C���v��`Hq�Tc���8 �)�g�����X;��)9��������YzRl4N�֜&���x�t���_'���X1�!�ϟ�5gn�io�,�M�c[&b2�O W�ݬ_4��k��7�';f�s}���a�o�>�b��l�dnAW��WW�||��n7֢W��&Y�7[D�\t,�lf����ڻߺUI�H_��	M����k��͍�M;�R'��x� eV<�S1�V�׺����amE��tc[=o3&�OMIA-�s�$��,�W���?�$B^��o�5�*XH������ ��3��w�C-2
j��r#]��s�0�W�m hX�	F�'�}�]�M��U$0`+�
���l`Ϧ�W؃�	�#r�&k��En����_5�yfr�xx��Y��n����Luq5Zol,-�L� ��m����)m%�KuH��6*[_U^�F�Ñ�c�ֈ����r��E�s��s�R`�緍<w_@��ًd08�5��sp�@�V�� �8@)5����m0&�wJ6��{#��\�o�/}����9�ڝ;��n�{o���U]���(��)�d_[�&�҂��/�o�a	�m�0<�8�#��z�Y&���xW�{�ޒ�k��A����ԑ���d���R�=�����/p!v0Z�`�`�AGH-_"��H\F�pF��3��Q��d��}�ë���E�3�z�����̉�i���O�����A7� qVT��*���h�;���71�a��u����.ͽ9]'X7.Ҩ�,�sԱ!�]b�f���`v՝��Y�;~����xK��;2�@Dݠ��"�ډ'�[�Gdg�9�5#�QwZ:����#	g@���S0c=p��ƥ =�/��0�I�]]�@�/l�5-�~-,������%=aD���>3}*�#&�YYp��������X��GA�š,�1<r��K�n~a_Ȧhk�q}P���a	�^|��,�;����	j4+6z�r�~:��FG����>����}����yI'�Ŭ����}�[�rJ��4�Z���$�%.7*��P�H(T�r9	�Y�-���p����L;�&�-Ҫ0�.�5����ͯ�P���,'�>/�Opx�uHj���r����9��Žgh�-��*G|�������Rr�w�+��ɉ�����)�?���]5�1�F(�(�Tg}�$��/>�7t�'dx�|�_f#��~��ԅp�M1�����d#+E�f(ӬG�;[�@��@+?9��!�j�6��J֪�9_\��4Vl�TM�!ٗ+�[(�� �< �$����� ���@�[�.�њe~��}-�O_�`�&iN�|��x���� �+S�M��<>ᚙ�J9iF�;YY���0�F�J��.�e�Ss�t�L`����D؆z:hp
qZ[�����Yr���)��d2XI�TI�I��8815ƓY 	 �d+� u6l����s��ޞl�������%�~������f�@�~BRD�xw�\g�/�g�u���CӪ��m?Ӑb�1X���R׾�ݍ��YؼD��8�N e�����wtu9�	!  �fzT�֢nܕ�b2�\܃�kNGB�������	qu|�� ���):�����I�yX�a�͹����_�D{x%7�pV�,G�� �O�f���JɁ�o72��(��?��#�{*\��ϏHICZ7a`r��D�%�.���I#&�5}AуGgv�<����އ~������e�a]J�f���n�E{߇*��׉���(�����Bm�m����:AXs( �9Gv�-6g���7���q&�u�E�CqWk��Z=�pz��B�CHO�*wCm�s7��Gpn"X�[�F5���[�-;����pF�e�%gU��g[c"J��������Z�;���]�YN`Xr��	�l�^h�p�pt�ԧ�o����	�js{��πY��).�u�zv�o��P�I�~��=m�o���4X�:�o�T�[��W�B��Z��LΚ�ha0PS�Rp�I��7bv
��5�ʿ�@p�� ��r"��C�1�$44�)�涷Մ�ov~�?񈊞����`��/��U.��Ȅ�--Y񻄍��I2+�{rGF�K�W�G|�8���E[%��s�%T�6�(r�賟9�,_F޸X��<ja\�Ҁ��h�T *��@	�em�q8ԁb
�/�$����2�ef�O�O�>���"|�~�(�M[��緐��f��3�M���d!3��_���ȾfԌL����2�ly7'���u��� ������*�����68k�Q��]/�)�1pW[�i�/��ʻ�?2:.]wV�:�Y��H N�b;��Fh�t�м��5F?ZC
�_j>��� �6|��	��s���̄�i�j*V��q�H�:ʝF�nY����<�����+?[�|Ej����~�7�9��ax&"��<���k&4��v�x�����dO115#"2bn�w��u �t����{��8��l���:�yU �z?p�#aa���(K R:�VtLA쮤8�p�4�q`�ܺDm����`������J*=�xx�=��>��t66���B�94��N����w�S&|�9Y�]%��;�˯%�})vd�#�v��^�#��"��G�߳7ۣ��u����>����v,�����'�4��8���o�~�Px�G;�F5�[�K����z���4�K��b�Qc�:v�`58��x�rU~G��g�҂qdw�Nm�A����qX"4��`�W�m��� 8 (+{�T�%���&24�L,�J�J*\l_.���c��k�ڇW�J���'v��n����9��wN'�.08�H������{� �c�j���JQ�����V�Δv%�	m��,�=v��u-�py͟��R��/f�1���-K��W�@�Q1���㯜���4e
�gE�3�f-u�:���d�vڡM�����Ґ)�#&,#`Xu(he�@�qV��9��*�f�������!�%��}�<�gr6�E���6WA$�0ʁ��d��j��Jʮwk�a����0a�1L~�\�����`��Q� ĲA�n���G�����<Bp5��H�H
	 �r��U�v�z��8X�h^�,�m9��U=Q�0�ae��!d.��-[����	P+m(��ƶh`J��i\��m�x��ro��f6+�����ٺ�?~���|� Ks$����l���t��HP���3ݝy��^o�x�v��ǧ5��Bo<��oJҗ����< N��V�{�-V�M�6����1�5}?��$��rҖ�-���<�S��ݦ�~x��j�#�;��p�i��z��|p����V����
?,���Ԍ�N8a���uQGXD�NB�[h�x��ҞMV(������iSC1ҹ�?9dG�b��Z^��Q�?=�#�p�3��ȓ)��r8zn���1:��������K��\�^�<����U��y  ����A��{-�h�D��/��̐ڱ�N�o����CpT�H��܎Ћ��>�/E^]ܭj����.��S�x}l����i.nfj��Z_��U�'e�~;�����T�#M���А� `��"�#����b�UI�%Õr��+D��V
�[�o�� %�}�F���ź�KIӘE�FHl8��g�Q�W���I6
�mtyNӃ=�������5j��7tt-0��d����)����L�p����Z+�B�.5h���oPz�Q�Ų!�FyJ��ɦp�긣��ET*����
u�z8�	��m�3��:V-Bq��'|��4���}��R��-��nA�|[�Sd+cZ�YR��T�rT��b[]��Z�BXo�2��>�#5�)��pV�;Qs�S��t�ZEia!�Um|��I���{�g[�b���Z��t9{cZ���"�a���Cс�	 ����L(*:֝˹�����^B)}�+�G,�������V��߁�5�s�h�٤���'��"Ŝ=p�FA\V��Xw�/��[е�m�S�.�r�����pARq^rG^$[p���
�c����EG�O'G~�����;���r���T]�M��K9�hǻ�-��z��k�Fhq�˨*����~�KJ���7�_����$�-�	�K��	�F� ���&�4���Q�҉�{��쎟B�� ��Y׊��R
�o�����3�缝�e�ٲa�c��r\�u>y��~�#��㛻b��X=�B�-hol�5�u$�1vh�۝�������o��vT�Δfj��*y��@{T5M�O�O�鯰�r7w�JN��1���Ek�E��쯽��+�[{��)��$��+����h������0�f��I{���:�^<�J��L�~�Z���G�����(:�(׻���9�6�a��T��+��]���hϠ,�{� �<�p9$�Dˡ!�pzE�b�S�����z�&^�8�����o��N���߿�"�m�g!pCH��C�"�����&ЕylF@���2"�	���վ�y��<�	Ġ�&�?�;�Tm��t��c�;-UES��K�&��8� �@�;��#�N'���}�"R��CKV���h�"�6�����a�N%d�\x~�6�#��^n�tpR�z`:�a�C���n��X����f��N+��д��0��̀�� t4�b��eW�(�h=h�+�iX�`$"<n��[r� ~��[�^��Z�I�+�1:�kV���B�0��e��·�n^m~&r�G���
֥Ner\�s�W��Dl�p�|�!�fp߬Iq�z���Iw��a�2�!д3=���� a=Q93�Z4'sA=�e��0܊i~���Ȥ����np[>�rK�����a�J��M�|R*�E`� ~�ia��Jg�h�.� {Op� HٗA��a�C6Y%�`z`Q>��8��MM/����t���˞1�͎�l��u��گD���AI����z:h�J@؝�]�z�*^8:%ā�*$�`QN�k�_v�Cgr�ï����٤��{�6w� W%�ڬ��?fΟ:x�g��mW?�r�qf�i���i����%:}���ѝ��(0Q:�_�6:���y�%���������(��|;oo˪�V
�����ϒ�T��M+ϷԛS̥CtCP���}sޚ������I*��nu8>轧�}���#�?pX� \@B:G��w�:Y4�[��d^o�U��Y?�7�����u���I���y��ݽW�}����e�)R\�ꌹ,�\��"|q��S"?4������ڡ_㪂E�	Ot%N�[�� ��$-�V���B��=���ia�<sDv���Q�G���� `^Q:�Z��Pa+8�0`S��R����
��UH%&cИ�f)�ɴj�j�u��̿�f��E$��끲��\s�X���x-A#ղ6�7���F8]S�DWHt�;�� �ս-nk�)�Ԝ~^��%b�/|�!�Rt��D|1AF�z�~����PE[kk>O���`���Ւ؊��(#��u�l��ӓ��z��;*��6�(��Q� \�nX�u=��E���PZ��U����$m8�:���-x~�<����w� �ASض��x,&����ـ`�>`�fp%/��\蘊Ԟ�V����F�|�@u�4�d58�Ô�g٨mc�o��e,G��L�u>��<��V�P����t�I��8"�U�wj=�k��&�i����\����O�s.=>�����G1�K��2�Dq\ė�2$bv���I��`5��*�'���:�:��L>�� @�L.�=�"��y�4["��O!s�|��'X�� �A3������p�m����Ī��U���/�?w���W�����r!��\�뼐�H<��@u���\�qa�iD̶ڡc&,my���A��}
]�kA"y�̴Y%Y� ��5'�`�
x.9���s4yK�P�����L���N_��J���w�n��K����:Q����?�jP���Ѧ窭�X�Mnk~^����?��������]#cgYT\,�Т����ѱ��y���+�w��Sy=W���^d/�����ۏ�'E�3�g�O3�S�|	�3Ϻ��,�5:V%x�2xS@��!p	9ص���1H �M�J���Pe̔�V�e�'�9��9�,,��AJ�v���&#3��Qjy�E_�Չ�2>���`�F�����} y\�X��f���g�)VH���B�;|�mVm����͝�&��SlRc02�ez���-�J�9Vv�x�P/���6�R7�=H��쌊�gS|ggZ)���׺oe���g���!i ep�<'�o��[ ��`�j8��X"j0�2�!5�,[l��DB��^�r����%X�6o̒����л�A�-�y������Y�|zK�_o.�p�Ư2��d넧;��W#����*�H�$��je�e߲m�\���ص7�nߠ�w���
`��tS�w����Eτ������5�b��
~�w��5�i���Űb2P�w4�e�F �O.��LX#���� ����������6<�L�
�ow,A��B�#4��4�� cш+*3b|��O�h�i����	����c���o'�L �׸�݁.!��
�ώ�'ľ��k+����	�R�)�HP�JD�=?����������K�O���T�f�w�0�[��}녎rK�m���ūJ�%��l����:.�Ɏ~�}<�S���z�r޴�v���@W'ix��v�.���{޵_nA_RӾ�W���Ɩ��&O�����{a轿��Ä8���3i<���]��me�>�pP�Kq">�y%���_����wy�L�8�{�:޹��yu�ۧb�#4�x)����� P�Q)��Y��w�7��]���[�H��+���z���);�Ԯ�̚�#����J�%Sԇ��W�[�x<$&�j�a��#䁑���h�v"1�sQ[d÷�PC�^�P�n�BX��X�!��:��h;K��'ѷ֠��=�=�7\���}��wƤ�{��ʞ�G}s�����б�g3tF�_�V¦CE�!�-��`.����|Ū��P��\����ʱ���ĺa�#e�Jɗ}2a�L0�[p��C�Fr3���}UNLb���Φ��IgGg=�>9m�1���IРϮա�XK�D}�^"�=L5h`���� biWOhG��U��զ$�נl���_�6���A>�Yu/u�ꠓ��l��t������#�j���0VE����u&0��37�#�����Y cC]�-����t�9�I����}���W2�6�KB\�I��}:��R䇛S�#6RO�m�<�4)\E���͔9����ȏ�k���]���k��m�S�A�X�e�=>u/ 5�ah�i^*eAy�b��Yq��Uڿ�|����%@s�lD������;4F [=����E�1Y����J|�M��gEv�N�]����/�x	:�����W�X4���q��n𿍝�����Ӕ��:U�o���t�a�����?���7y�B��L�����I̢��]�q75s��X ���/��_O� �{M�Th��?�n�ݘ�߇�Od�z�_��-���7�b�H�� 0��=����i+x
�d����m$�aیe��hN:�H�h)��+��ʪt���ğ�fIȷo�ˤ�e����5�Պ6x��g�O�	&���V�;QM4�99
̨�Ϋ؈80c�.�U&Zt�wm�������;�bNJ!����f��Դ�� B�d��KD4�>�/١Z�*` X.Wզ�S��Ͼ�Xŉ,��i�a> �|.͹���ְ����Qʯ��,����+��gF��G��9Vb����e]&RY+l�<~CB�+bݮ�'���nǙ��ř�g�{�h��%"�&���\[J����I���.�D�M�gJ�IDৎ�L�"�G&��8B��-��\�P��b@S�.`wӊ�D�&�KHõ!%�ن]�*�c�����'-�lu+bww�E��U�V�!�-�A�EW"��&?{�x����Ռ	j�h�h���+���'$�F�r�QB+#�X���'@w����;�}w�6Afx�$��]8YY�a��QO�����P,vw�l�.�9R�b7'��K���Ӟ{���V�E�4�@� O����4=��3��)|��#O��cNN�-�"�fi9p�}b�>�i�y�g!�%�(|����3���=Z��ƥh��&�ɑ�.+KZߋ���
q��|���D���2�h"�ӣ{�_��F�~�����S0����<(S [a+%�����2��U�z�I���`�X�G�� ���1�:��L�\��^��>J	-@�i�
�U2_��y_٦�˚K� :���&)�J���������I��#:ԯۚ��>4����{F�Wm�?@�A�g��w��@+83E�Ɗ�0�&n�gG���	���6Vf�_��c�;��ho�T�Y���=t�z�ӡ���P�*��Ç1�Y|������)���T��,�-���F��͠�R�E��)+�D��x�*��}�v�|ߞU��\=�)���yÎ�w��k�{G��9N����6?����v�Q���AA���,�:�NB���,�L�]Pؘmg��4���TP�yc`?h�#e2��DS�r?��<�N�F�t���F-�:(��� u�t��jKT�����vw<s��/��߻�"��|���}��� ��҇�@/Q�9�3���z��P*� �ݧ�-�d��P�Z��a�R�])��0�}|��K�����H	��ƿu��<D6#~��*���#��Ū���
z�������R#u������^��LC#�U�S����~�����l��N!��Y�~x��>�Va_baa�?H��s��ǳccV�ЅȣǞ䩠{w���'��>܀#:�6��m��%�QS������[&Q�%��W�"�y�y��a��=T©�ѩ�`�e5X'���$� �>��Fq���0�ҳ�"op��58`��������*��2����Q�N=����t7	���\Ao��Q�
�(қ2�}	�"#oD6�_1,(���0Nv�� }=B[{��x,n�fb@JJxcn�m�ݰ�SG�f]A�g�E*�=����������p҈䵞��� L�+
A��L:�t�)��8e�B�� (��]fg��}�̔�hfzEmFuy��6�Ve�R�_1�,��OSsj�a�@lՇ,�o�5�g��S9kڂ]Y��0��B����X�>>�^��w�I����oJY�*�����6����N_�e��y޺��En�-��r>����n���̖E����U�D�w_��D�P|o� _D�nh_��y|���<5�Ji������!�7t-_O;;�e5(�@_�>���J�|����% � :��.�8M@�\��"������ja,���ڄ�����vT�*��&��o*�_�Mi����w���6�����^�q4`���"t?�b�<�ã u�m:��:�ѓT�T ��`�x����vv4;A_�}vSؿ�6�\\�%7��s��>Wr}1L�i�E�����&�ȍ�X�Е+��;�ƍa�ݧWԏ�*mh�UR��܍+~���%b�9�Ҥ�<���,�����T��,ZcuP���"ľގcO?����]�=�b��^pՆ�뿮���Wt4�Ns	�Q{T��?{e'U�H^��t`2��{��r�����fzT���D��hUm���3`i��jQ�v7����|��U��~_�� �y�������Xգ �;����s4 �k��⥄����������ӈ��ٴ��%z�4�Et��7l�O��p�n]bw�g��;_eMy�Ţ�9R��?l�Y|3i$ϝ1�.��r��q�4m�[�ʅ�����	��>xʁ�2��jo�X	��Ӻ�>)���P*���?53)���}FY�<�@��G��BF�s�p9����:d��1�[%�P[F��X��-��ך���C�uX���Ml�/�m�"BC�9�@��Yɒ aLO����E�R���}�HZ��?t�r��({2�y��\T�������� m_���q���}@����&=���Wk��2\Mަ���㓏'a�� [�=��[���;s��m��Ҵ���*p��s��a/S/<����B\��q:3��aMk���VVou���m½RB%���E�N��Å�>K,�Z%z�P���/���x(�����<k�};/�p���N�&�����*4,
���Ac$+f�5)�YG�Pn[�J2��t�F���A����6'�S��6���.���j�j܈IG�3���ʒ��Enc��Ot�gC~J���~.|���Np��C$�(��nG�0������u9ši
�.��my���u5yO��2������rul�,&���:�1uI�x���H�j�8J�붆6����Z`P��Af_Xr���98]U$�����o�`x:{�a���9C� �n��?T�iD�s�fʓ��!��yd��H7O�[e(������H>Հ�:�=mb��>s%ry��qݣna8$`��"MN~
'�tx��k"$Ǎ�x�n��8�E4�E?;<�s���&�p���E�0���='�η@��lH`��nn���E򪭗To6^����(������*��Kه{M9�Q%q�ȼ@���9��뀣[H��/]Í �{o�(�60F�w�0S������ㅦ�͑�W��i�gI�E�p�n��yA_K� �-��xW=�3��^�J^���R!#�\���R;����0�������"�H�g�B4�{�۳{��䢠q��E��8�E�cML���-s��6����~�2v��OWs<�ߨ������e�0����JH��5Ra���՚:�g��3��m���t)d�f���2'�����8W� {,� HH�`�̬��l��α�!W7n(7U�Z���L1<P�#�V��v�Y��e�e9<�j�^��A���y�B6��t6�E��
�R=#���1��;��o���3�"Iwh!V�}���_��x�C�q�m�Ex�p����#9`�.��"��F�`��?L����X�θ2MY<F/D�o�>���1��1���t1�����>�m����q��%\.����(�f��N�₆���~��ܦ�I" '�a��W�k��	iO4����3Q(@�	{ݼ4�el���c�ܦ� ��^w����[�ȕ�yZ���w�	���HԴ(���Iu�	NI*I�
PZo�R]kub�)W|f@с̉O�MTQ��%�s�ʇ�[ޫY�m3�Ŝ¤\��	����l��<����7�Yy:������j�N��~�ӓ�͵4	���C�8y����$�����;�����A��=�����ōx?���=����-����du�X�B�y����?֪&�=nӺm������f��_��M5�A��]P��~�A��G��%[]��Hi.yq���%�"��ȷТ� �;f��^��c�U+y13�_���5Ƽ��*���Z��V�,��a5�K
N�<��Vӎ5�7^�HWG&���>�%F���� �~J�f�wyP�!� B���R�H����]�taRF\�+w6`ఊh��໨yI��T��ZѬ�� ǘ��\j�.7xD\:srK��	X"x#�Bs?"*�x��.b�6Z�r�Oc�sD%#i�	������'^�t��xQC�B2	��x����%VD�Ab��X{p�L���Ԕ�R6ױa��.dvےChLj`��҅AR^QRi����p)\ό�9U����u	���G�����u�s&�lq�� qf*	(1w�pJ����!�M��T�$�~j�f8���T���Xc�hƢ���f�w{hڐs��1��OR)g
�Z��-�i.�u���$"�yS��Ɛ@�_�H�ŞnS�ƄB�&�c�f���2�r`qʍ��/�����?�v��Eh��C<u����a��Quv�݉KL����Z��a��P�M��!E����>��.K$ծ�F.o0�b59x�]�H�n�mb{H�1���<]�r�0�K��"�v�Mt�w߼���������2 �q^VO2ҍ�RƧ�������7K�|_t�{�#����!Ԃ��c�����.�4W�:� ��� 9��N�Ձr+]*N��yri��
N�:��Qq#
.$�ᝍ�Nή,Yd�E�g�!���=�Pq�K1=�ti�6��熀H���0֥��$��C��"������K�/�RO� S@��(f�  K��Dx�c�z}=\����4��5Y��T#�F3Y�mbb,ͨc������z:	d�jמw��,���Y	��6�P8��ѣ���r�AN��Bw9�H$�GH�z�m���tH����U�A�η���0&�r��o�%M؟��v�"�]sܲ�C�U&3��pcl��h�	W�(�7�K����&�200�p*�Z~e͘Ac�����ᜑ}�C~�%B��x���ԫyu��Y�S�Sa���ܪ���s'P��s!�mU��^�:���J�v�@�چ��i���z�D{~��P�pC ���Ȓ��P?�PZ����q�B���*�m�4���;U�Ǌ����i�V�5M�ѽ����T���,S��ړp�ٹȿ��f��=ը����DZ;or$}��w����w@�e��X �+�P�_�L�Y���+8������xm+���N���i�/�95��1rM�?:$˖�T��d�B�L��r-@k�t-[n���lZ3v�g5�����S�K�յ�N��险����ޡ	5#�fM�*�J�����( ��Yp����rlr&T~����<?2r�}ݏ^�xq�f}s���Ң����*�cv��N��� �.��,C�è@�~��p,d�_���]x#��h�~[T�u�^e�iq�h��߀@���u�B�k�� ����Ј��P9�)�	rV�λ�>���V��'}�W����?:2(���C��|.�x�7���&c�v�õYH����������5�t&�҇m�&7�ň'*�*�eD�,�ދ�.9�wp�^U�]I��K�����NˋjN9�������6�@ ��c��m��i���|+В�]�������8�z�f��(��6�1+�C��y������ߟ���C�����'�H��$�C��q!L��,ʹ�Y�FtU-���F�#�2y�sv��KAtiw�L��_�Y�b��^9����[oQ��D�r��Zt4wk�b h�u�ޭ
{b�e����#|^�du:7�r�P���DZ��n��GߠAH�ѪHa�����r��Ar�Tk�� i� �a5� �����|.�Y��Ω�=���n��~@����N��z\�]_\�ɛ(Z_��:p���۰(åX���sY�9ׇَwC��L��c��%���b����W���hֵ/�յO��~d������1�<׷�s��=�z1N�ғ��v�@�m�-�����},��{���O��º��}Wf��Xo�L ^h_Ϯ��4���s�yW�"�[�L:�	�9V	D�zq���P����1	�\/�����b�R�"'>15�z� ����T��jǟE��.9	�I["H����Vw��hw��pв*4�oϔٛP:�o�.K=��'�45H�r�mT�柛���ƉT�"\���S�Q,�e���9��M�U#�oʎ!���f�&#�0�Y{g찋��i���@�89�A���"	��?�7�0'r��5�������?zq!@m  �}�4�<����`@D��@�;��1kC���*T3�����&�mM�����n����i*6�ؽz�r��_���#��kf-ֱ�P��]L�l�0#S��j�:屶&�b��bB��:�p��F� 5�	�Ҭ��B��Ƚ[k�(`,�?�b�:	Vaaw<�X�pS�ʕ+�6B30ҳ��=��VK���P��>��';�>�E���5+cg�/b{��͘t�^�0@��2Qf��2��Y�u3[Uؒ���z�h��@�Z>�ܞV7��\���j��\���s��0\�Cc�5�����n!Lυ@+�m�\����U9��aO��(u���՛��{���=ۤ/�m�>{���_zq��K/�Mm�h�L�.���z�X��l��-L������j-�'u:V����ӭ��_��{WG��e��~��?�Ý��;��TU;A�/�tҋX��J,�츜�~TP�M��U/��)�[4�Wǡ�!Y>A�G�u(�ߨ���3��(�	2(ǍC�R婢���K�+,A	'�~$g�Q1w]z�^5b�)6�֌��6}�\_D��{����f]ןw�8	��.��o�-k���t���erh�����{�a�����]�=�`"���&��Qˇ�~59�m��^��^��q�+X�b���]u�˖BP����+$F�*���rzw�5�TO�j��M��O�]]CS�!�CLL���$}�n�Nni��E�D�[*��8�l��b0N�)f���U]v`���垚��r0�%���p�  ��D�f(��55�%X�}�ݪ�/���ZS
:�������ޥ�9ұ=��ݸ���q��Ņ5��ID���ؼB�#*2����#mN�7�X�� � \4��u�o���I[CM(l��q��CwܕF����}�u��m��H[lS�&��� �ꚇ<���Y��;������
�T0Gp��/τ�JЇk��r�M���.Sf��6�eKI�E�"2�2����yפq:��"���E�G
��U$���� O���"�2�X#��B��&�� �8/�H���4X�@-q�_�T�0�f9�V��>�������y�_�:?w�ڣ�;4�e2�:������0s��_I�ź�����3g���0�,.��'����/������ps[ Vs�[e ȵЦ�ǩ��&(LЍ��u��U_]�O'���ban���������g?����c7r�����]��Թw/�5ok*'��:&�H� 9�S�"_�|9֮��� ��4v��K�8��[��k�s��N����#���ɓ/{���$�fG/���Y2��$?�����̅��y��|��y���P	N�U
�J���CӢ���4 �;�c9x M��h��.u*X�����Ԃ�2iP��W�ޫU��|�L���0��昄���l��$�rS��v�B�����#�0���� ��Ҳ �A����-���u�;k�K�1��$tI���!�z)]ʘ�����nyt
�9�L1ދ��ՋWg5�,�œ��)�4�m�&�i���t���������o	��)8Y]�0[�*$o]�����{�ź !!%eb�-}]ʺ@цlD���	���3_�~�$ӏ!<q_�i���U6�@Gd�����
$ˁo�n���<���V�}m�?�oJ��U���䁽itp�
�z��#[e�86D(�ׇ���.g��8���� X:69�����!etNkP�bΰ��E�%���
@�FL��h�S�Q��� (��)+��	��gY���@� ֊���	�~���`.�a�x��t-�eNzl�NԵj���_�X��?�A��g����kg�"l�ư ��F�p��E둕�F�qr�S�\^��xy����:�Ǜ������������z}��ɩ+��4�.Y�@/�����@a�nd�叚͍���b�=u*mJq��c���w��#���{��������;�n(���O<��W��b�����C';�X�X�^�ƭ��nPQ�ОR��5����bi�r���e��t{��(r�+�)m5P��9[M�1��@&��z��!-^�@�i˰ �p��Y�s:.ՙf`��5��w�x/K�;��g��t%�hGw��A�C�R��,J0��z��l3��;\-��_W���.���~���߭��}��w��������+W�SC�oH�N�11H�qc\u?_S(�P	!:�X-9�����ѯ� � �J�d��^ W��e�^98��'�BtU�!�\��ظ������L�;���W%�S �*@�B��M9����@�K����I4����q��i~v�z)@��� ���Rd|�7WР�+ԴSW�M�]�{t��]�>7�l1�tbTsDc֣�u�&�X��\Xн"�G�Y�B�=
��Vaϡ)�ɗ�m��uX-1B0*�T�]ieiũ�| Ƹ��<�P�H�����s�q��=ڠ��F�2G�N�2����;J7F�u��X^ﳸ���H����c3Y�q�@�!Tيg�Ws�pd��fͤ�1�d�i�gf��?l�� ����s�'�rdm�g��ҳq�`��
��0e.x���v]a���J��Ԭ[S���M�c���~Td��̘7Ed�a����kЦR���
k���^�xׅ���Пnh�l��������կ���wv�ٿ�MBؗgW��mnJ<�F��[��Ȁ�[[���fkx���v�|:����8r������|�Y��çV~������K��S����������Y��U �充��_��^}3	��3��עm];�*��~fg�BN�M6�������,���Ԧ�yuo�������a�e���9��ےC��E��\#���+���8��a�[�����Ph(a
�[�.��|�t���t���ZT�;9Mv��zۡ�q�P�$lA�X��H%g�L�$r-�-�{U }E?a,]�>90 �-��:.ߛ	r�O�&��� ��J�._��hٙZ�匨��y��ŕ�:Ir�j�*� Xrw�B:h|�1��:9��uσ�L��{o�����43;�ώ��4oս��3���t�%靖�c�СC�J
�ș^�$�K�s�2�]^Msr�;	-Q���uC�c"����0R��u��J-=�ȣ֌�`�ˈtS[�FM4�!�]��bb�����!����T��.�mb`� պX%��M�T�����S{(�B���u�8ӼsQ ��f0]�z���u�
ѷ@���eؒG�!B�U�	ז�(��G�L�u�G/��@����C,��h�4�7U��9�s���4{��_'9Aǆ��x�N��F��:��C�/����#����t��c,xh\BA�D�i�����8�`#�fԵb�<ﳚ���]�_p��!9���-6O��ļnT,������H��F_X"�%�7`��`S%$��o�N�(h�����ϼtjߛ	�}��M��߰�1t`�>���Ƴ.�*Ҫ�R�gYi�P>�{k��nľf%j������zm�t[k[�\��z��z�:z��ܥ�?�����W_|���/����c/����=�5Ϝ��]�+��.IMH,�ey��A��0�p�+v�!y�n��&�푢�ȱ*��{��5��%@�KA7�;����.��pMN�`Y5 !�
A�5��QU�M1D�[q��) <��������9B\�1q�d�hX�1��O�:)Ჾ?}�Y4���1�(��% ��sx7�Ε,)�'v��!2��˸Z����juP�g?���H��+�p�E!��PKH`gPi��r7$�~��w�xG��G?am����L���A`}��ƦT�&�%9ܤ{��Y���k����>1}n^sO������
48�k�SH�G@qU�G�����2Kb�����ۗ����3��+�=�t�ݪ��e���#��cD�C>8��b'fu{U�0 �yhj�$2�z �-�E�ی <x�kl{)��sN��7���-�m�2�p��b}:� �T	�����vauU�"}��`"�ȨD�>"�&Р� ���+��d��F�a�*��ӛ 0a47�uȁ:�0��6�Tz�/ ǈ  ���Q5���`�(��ЗXBh�� N4i�/�{��y�#,u���͓Mh�gw�و��� U�
GP���:��<+;
�}�a�^�f\[X`�8�`������*$�s:�ԋ�.�����9�������S����m�{��w���/_��n]�ҕ���ͳ��_����^n�ru}���nÊ|m�(���
����\�E���( ��Ya�����`s��ٱ)�ܯm�v����ty���qG{��]_�¥��w^ݜy���w���G�?�y�܅����/�����R���I�������{�7�Kޗ�A��! i�Ԃ(�Eتg�H�4� I~/�6�P���}n��Խ�&�8]vt .^���6��FM٧��V 28#��������3�Q��R��Q0�U�Ē(\��eP�s\�����k!ޯ:;_���Sȭ�Μ9��^�p�@�;W��v�G����c���n�W[���c��iF�߄�6u~��%�!?|?�,5v��ջ�p�k�ȹYD�#T�lU ����4AZ���mͫ�Z� ��_[�2��Z ��x��쓘�k�:0b:>E
�)`�莾����*���9T0׻���m��B���o�٫�g��x�,Հسř�tE 
!�18�3�O�����I�ti �^a���؉q���Z��I}��3�
p
��oِ&��~t��I�L�&���� ���d�l�<=����Q�n��,�� u�4�\t�&�)`��qm6�O�1���4(0D�!�!�nB�͜D<LY�Ua�k���)�Ɵ��^Ը2["�d���˳�>���^��#�/ؾi��\HT���	����*i@S{��ƭfh�C��٭B�yJ�g�}�-/�EU�� |�wb�`�)�1��B?_ ��B�CH-�������[q�g�o���k䦘�Im>�?�*���}� qQ˥3xv	��xΜ�|�	��LP~���H0�`���b
�CO�r�;�xF�p� ����Ͼx��l���t�*KG�i]͎U#hKu�J8���[����i�Z]Z�������DOtO8�٥i튺����~�l�볏�|�q��~�ѳ������_fYZZZuy��ѡօK���]��/<{��^���/��k}w�M��C�.�q}�&C�#9;z9�G综��"�[ٕݫ���� zQe�@���ȠK��H��%���[HѸ��DÄ�/�n�]���^9]8%�';J�"Z�I9:�t�v�rh}��~#��! ��}"�$J���/�O�iT���H�Z��HM����U-�����^�i��q�)�%�)�(����n�����{t��n�)]���0�ːj�cg�V��|I iXί��7Ȁ�C�+#j�H��>�����Ki��ai�4
`Ɏ���}���<k [r��REZ��@sd�Bx.�h1�@Oy2�hbz���� ��YW������[�#%d��Vh��2� Y�
�"<�S���� �`�cj"t@-R��rB�~疛oI/>�\:������ �/;���Y6�FTǘQH��a�%�f,cM�l
1�j,�լh6$���x�)(�j��a���-
X�	�.�C�HE&]�lb�r������ƻ쬪�{�S�R�{����u85^ǣ��xW�I ���B��7tx�kI�^P\���� �M�W}ֆ$PG4Ӧ�C��l��#G��e������GR?�TU�1��EB�+��f���8�D�+�a����P���0�{��E���[@v�,�̋�Cb 8�72��[�!<��<4E����9B�6���nȎc#���S�>�G��~~�G���/�n��Ͻtf�?|�_s���w5}��m���'���P��(��߭�߂�+ ���Rc��T��K쌲�Y��ؐvt�[Z��n�觟�˟�L��mǧ�>�w�5�SF����։ڶ��陹��/^�������zsO�k|O��d���� ��j��UP�r��71��U��k!�p
y��f�m+䑛��Fm/�G�&�jȚ{
qy�J���q�uQ��.b)�ʢ��ށ@uJ hM�A�4���ё|���8~v�%4h��uEQ���Y��an�Vt�9�1�o��Κ�rD�����m��:<!G?R�3꠷������i��&�_�u�`�E8eP4�ژ��E��;8��r> �6a�q��M�kn��F�K�c7�<S;�P�����*��4.���^��ka�t�ԅꧾJ�o	��6:1�9��0�Ì:/����(dCas Nw'�;1!�e�\������c0 [b��*7�`�j��1,ئ܂�Ԑ�9wu�B��������P%����!L �J����K�|"s�7��8�2<O�c�l�y4�7sbì��h�^��,ӳAq�,%�ܚ��{�
����*�H^�bUz�74n��1�j�W��P���~O�<�8�p�N�����s�Ⱥ9�j�*���bߩ�f}U�D�N��c��}�{ҧ��P����κ���[N����t��e�ߓRާ9�����s�L(�[�d��q��% hvthɠrU��}#��w��Uq~}ܫ�C1ǝ$;�ݐV��. ��y�r����[Ͳ���	�[-(F+��C����ە�^���0SS�T�y���g���_���+������B��S_8���#z╙?��8ᢝ�h�	�������S)�Kw���z�X���j��;;]���E��F�9��ӶfqqV@H����������j/��Т��Š)jޑ����-��Ԋ��58���%� �j
���&��P��m��HD&)�A��a��Uy[���k�%��r���&rm���Br���h�A��� �ɉP���n�2T��Q��sreI�Bv�#�ͦBAJ�v�m�1�PMyU}���Qe�W`lP����)M�:��!���p=rN�>�.��e8s	8ӱ"<"����@�uK��#��R�ՄuPE�n�*F�������j�s�V�, �F
��a�
 ���X$ݶa�1���k�JӃ�"����;�Cwݞ�z� �<�=�E�V8X�`n�0;�����#P����f�r�NQ4��!c�0����Q[F�l��d¹Ѯ��R��[�@86:��t�����{��w���S< 7bu�"3��[�ǚ�քlҒ�V�E���b!��B��v0Sݺ~����=W�/���s�p��!�?SefFsJ��� ���M���t��8;K?��ֶ��*L8�1fR�Uf����0�!�ߖ>��f
O�H�����mVl�����
��N����4���.��l��i:ΨB�\�^�fk��!��C��u{�G���{�������<�������r9Z���|�'���`\� �>����P�wܮ�E+��f�B\<����d��b�=�^��YQ���@�l�Z�3N�s��f��0&`��lP�/��4F�W��'^�x�;��~}�G�#��?�'��f���o26�?�4��ǟ8�����詗�}{mp�N�bִP�����G���Z�y6ހw(}�X���)�5��r��[E���%�a��K�,!#i�H	��V=.4yZ���%���$,�&���f!�3�����"�ϩK�{ׄ͟7�;l��D%H�LU��͒��0 �M-��*T�ӭ����N�u��3`$X>��I��#�MιWkLNAj�H�k�f�,�d=ձw���a�v�vؤ6k���ظ���`���B`4 �F�@�M���h���qU��-��5���V5"�W$2ݡB0�b�&��BK�8i���8�
68�jEa4(�=����)��J��nK���+M˖2�`H�����G�gj<�똿��O؉q��xU��;�X�ʳ��a��L�
�-�w�
K�J�C!T��p���7t.����W%�������0g�*���T��R�]�>X��]>sN�D��N�c��)|6�N�>�fp����P7�y����׮^1���1H :a:�������b� �d�g:5?��F�
MY5�PtR$����p��;��M�kM�)�Z��6�j��{*+S�ѷ~٥q#��0#�6��'�ӽ^R��3ʜ���U"aX�V�X>3$ 5,�CB���Çһ��٧n�'MپG�}Rs����<M����o�`���H�H��]ߕ�x���_��N�Ȟ{4������\���10�^/`��/� �� �Z��n�� �C��Ue�e�b]���C'hh�z�^O�iM�D�
�D�z�y(|i�yLs]2�pK]$�<�~q�q��*H �������\���c7]��<���w?����}�C���=~�������Z��v}�5;7ףJ��Y�/mn���|���ϝ���k���&w��u��7��Hg�iS��R��Em^Ƈ`E��z��|���
����I�qy�v�n���3�I��V]��V��P���������ve��q �}����M����dQVl��4����ܪ	!�v{<�tp{R�go���oC]cqvb�@�5�aW�_�>f͌Ő,|�k�R���?�A��{�43��F�ێ�:;��SS|8�G��h;�$T��}����#��	-�	c�1��)��1��BȶbJH;v�\��y]�������_\�ty	R)�뱨[�G��'G�PkR�	��F���!�#骄��W�l�!՟+�r���v����ߚ&GG������@�,�ft\ q�@Ì����u1(4UȆ�
C�B!AtXb>.���Zz�q�'����!������ 4E�CU 0���uT������ �#��"m�����(Ao����F1r+��G��Se����6��/=�������'���~���/������c4�� ���#K0|&e�kT7�J̰_[�W��E9�TB��}6"TC��ǳ��>KU��Й75=#�<0O��L뺄�u�fkn�q�m��<d/ ܟּb<�~ �s
�ql@���SW�?��e���GD�K���ӫ
�1v�.�"S�Mڿ@1��*[����;��/��/x��]<{&=~<�sN��tt�y�7��Ok���ؕP+��
�m�؆ ���d�w�D3Ã5`-yV*@��5<���E?<�4�!�}kg������f��3�C������F=У��Aj]`N��P���t�ۆ6?C�#i�������S_x���/���-�/��412tq��{Y�9����_�z'ֶ���Ӂ���}�jh���z���#�$�k�	mh�ԡ���D�ʁpP���&( �Zi���ROR�OU���kI��שJwۢ|����C8��5i"�{G;"��m����+���C�Bq((*����wMo����r�G2
���
���o��D;��r-��a�X��q��íBYd-���m�[8M�O|��r�E;W��]� ��)8�7��ǽ��̈́$h�J�⊲�S����a@��~-R�?�,�*2']��3�tk��.**6��!W!�>��7xw��w��ܣ�e>|"���:k���+N�)$��g`�X|7$&}��5�4�b!	�j��.!�gD��ij��E�����+ 37�=w:���}����dﺄϑ^/!��:�ώ����ү�c8ɵ�p��38vv�%�Q�6$�: F�R���z\����)a=L#U�	˸E���w�}Pņ ���MM-a�:���/_��&�����ߚV�i��x<}�[ά;�����C�/�ȏ�����#?����F�3?�����E�#G���cH�N�-8�m�7Y�{�x��x���"�QsDv�w���;xPUR��v��_`��KEl�w� @U���_��@}v��"g����qL��[��[�G>��Qi�n��v���<ux[����fc,u�[�X��皀Q��306�Ω8�ɓ'U�aX!�=b�V�z@�$�x�4���j�K�ږt�9����b%���P��N�E]T���$JB,�� ����#�N�R��Q`���j����5�c����F�����
��i-���Xd͹w��+�Ω�Lm%�{t,6	�kZ'���|���0�59�n�=�|�Qe?^M���B����g��B�H `e_X#4}5٤wd�Ca�	i�&^��|�٫˭������JmyeY����>mV$$�JkN$jt�Q�:��^'ew�?��zV�=�hú(OZ^ot#͂е���"ւc$�H�|l��x�q�#W�_�B3�3���C�(Zv����{U�3���K����U-�v��?{{#��k�v�.MO�X	=��}��4,r�Ҥ� �]8Q� �%V�N�]ZP��H�eEK�jA�#�\���fP\0�q��:� �/����pֺ��%���Dz4U������^�h9��JA�-?f���%'ֽ�/�(|�0v@�uZ�F���������4������+�@v���e�N�;�I��.9����O_xQѓ�%���чK�+�k*[`��x��=���`�	�jQ��`�l] �
��(T�ۨ�6�����)���q�Ua��0�d[�Z�7&a��b�L������.�z���~]3�$�x�%���]L5Zq��E�� �%��:9�}�t�=b�v��4�THqD�[N=�E�tB�k���Ŵg`8���黾�}� ��!]�~?�J�����k�腆^��6#�J���6��e�>��O�6�L�qe���Z?�����eS�aCs�2�C�أp4Yd[ꃖ�����:�������O�TZ@޻oOz�;H�z���=\!m>�˦�����Q���i�� �L�Z�RqC2g��Tl�@tՇbp�;�p�E�n[s�3�(���X��e�>U����U��=`ʤ��D��}#iVlO��-�-�_�L�{�i.~���(ݕ~��~>�]��z�[��a�UϘ#�$5T���Yj��㽺�a*u˾+*�@B����J����P@����г��u��1Ӝ��<E碤�;v�q�7�<���s 3��\e7j?����M�r[4����ξ��eK!C4H	81���X��.k��jy��e38D�����w+���
���fCыSr'��@� +��C>G�H�"!��}����^��ya����L���E��>UhF�H� ��P�충�B��.�DMi���E�"�#�^;n QU�gE�2炄�iȜ�E�:�j�ǖ���X������g�B��ٖSǗ�P�`p&�ۡ�{�q�B �b���Ҏ[�ƃ�ɠ01���؀��%�h�9%V�N�^ՠ�Q��bǉ����t;r,��K��{����Mkr@�I��U��Bs�!<�0r4��I��~{�h��-?ܣ�
b�X!&uF֍4m��uL
�c<�w3U���3��y'��svZ7�
 �<R�`���&�T�|���E��c�P� W��a.IɆ��r//9�m�GCW�W��2FT$tb�;]Z��{�x�B�b�ݿ��i�����8�#��7Zp�۟hr�O����������N�jc
�mi<z�:�g�L���!�	l��k,��@8�K�<�P*Y}.PIͪN�	1v8{ݛ��%�:>�%��M y�,p<59��7�g>���#{'�J�2�X�M�f�3�M��9��@V U��}�7ڒݩ15,�熼0pKR�́/Bl��X�O�n��MR��w]����V��l�;�i��P�ĸ�i��yN/��y~/S� �K���w��xK��ŕF����*}�S�R�	���)h�A��c]``�& Ê�:F�\x]@�j
�\��i��g_Nt�Kk�N�"��=�&[�����7?���g�b�ٺ�P����s9��W26v��
c���ye�:�#z��n�_�k��$����d��i�ƌ���
�Q�b�����釼	����|��b��nl�x��2����??���y�����o�V�����{/ �;_-��Z��+����E�aBX�nm�`�i)��8�/g��"�$c��=j!�p���.�n�m�(bs�WHyMC8?t1>����]�'��ӭ�#������I��c����Uw�!jȁEJ>�M����)�]� �4�u}�
S���܄ T���rP��#
mP�fa���Y38�#���gt@0`��I�p:q�z5���w��G����\Y��i1�7���P��>ir�q�r�b�?�}������,ׄ�c  ����\ǖ��9u�:��}�^��Ħ]�9��Y�#��#�˂e��|~Ga&*�l�س3-\&4�ݵƆ������bm����;Q&d�x�b���>�������7�QZYh.�Kߠ��(g�/�G7�����t*�l2j!Q`@� Ӳ�#��S��^B[:6��v���(j���&�F�} f4w�/%��w�l:]���ۤ� R�歃�w���0c��������A�Ic@}*� �0�#mK�#ѿ ���u�z���N�G����QL���^�/��M�$<�-����Fu\���U���316,����;��)����lBD�����tTz��Ӣ����?�>�ɏ��S	
6�\�L��B�� �QK	^�ƽM�'�L ��Xy�����+:<�]
�څo��*9����VʆjfQ���t�ٞ�^?�̎����Y��τ�d�pi^*ɀ���b����#�5Bˇ�lS5t���P8���Z��	������[��`��nly�ՒC�a�[���A���f���倝׻��R<�;Y�p�|�ز[N�L"hkJ��f��7��� S��K���X�U�5�q��r�0Idn�c�y{���GU�%~X���-��8�馐��:ęjERA_ b��� d����s��zA>x���Y̨��ҏ�M��z;UdN�	���X����A��eǣ��K���R}���p�8�9���hx\���k�I�%ݚݤ[�Ȧ��I��9��֨�ZOVZ��Bf�<�v�q?ts�4��l�����y���i��ElN���zE�����ލ��Y�T���@`ѕ�->W�E4%�#(<�����;��u����l���q����9�9����	4�]��;��[bs@eS
����%6^iu��#!��N��^�@�}[ N)����]I��@ˉ	[��iga�,���$���c�-��"��P�pC�7�
0�!�o����fz�;ߙ^y�e^��, Y�g��S8x~i͟!�kR�9��4f�}��J�M'z&X3�l�
�~�7ؕ��W�Ƚ����k%T��.y��h��j������[k�n�1D�E���*�`K �B���*�wHn�>{D���[
�1v��`t�[b~�._��a�nI`�{c�cG��(��x��q;�*����|�Nic0�q �![�HO�K	�I�@�'p��Jr����*�S�T��:6��C]A�Va�j��F�.�X6a~����:���g�}�h[!8��"zD@�((�c�JB���ࣜ>�ETscΡ|��a��n`�x�[��(	-tR��H��ubb�U&^���o��Ui�o�_����@�Y9Z�W� ��	ƁE}YRT��U�R]�(�n#O��$h.efh׫�&�+2��1�|�j����S�0 IH���/�,�\C�
�[ab�u#J��AP��Y_	�H\�
��n \�cO�p_C�+�{�= �Hq�����PX�;�M*���ZG�Цt���Bg~��qũ��Td��g����0 �r�M5�DD�����Q�ٴ*��C�K�(Ш
F��@�)�+�}c]�D�;�ޏ`�����j��F��p�a��ơ.P�!;8=Z�min5��� ݒ��k��Xֽ����n�д���f���}�I��ݷBH�
ڮ/�����~^�O>��3lV6�R��tVs�c�=�
��J˲��y	ʛ��(F��9���ngGV�;�H�B����s-Oy�7rO��+��ԔTP�¬�����9�9�p!��t�^��9��QAS��W��{������v��X-TY\ ���KU�E���k4��(��(H�z�'m��XƁ}ҙgt-l(�R�#��F��~�S�%����Q��4x��y���[o�5�^�v�i�y}?41(���A�*�y�D�$-�E��F4�������WU-}%�}�-�c?�yN "|�%@��z�E�hj�Q������2u�^(e����j[�c��L�U�9��u��Ɲf����Dk8�B5�X'�>�M���r]2�����~2�i�b�Cm)�3F�\N�Gn��9����,�fэ��.��_��\����r( ��L���'�;';0����:���[9735~h_���9u4�Ĺ�|8��_�f�����I�����d1h�;|X��g��q	)������i����y2�^:yF�W#�w��2rX(�q�,��	���>-p�C� U@����&V$�)�J"v߱������\�h$�T]9���hT4Qѝ���v�P�M�����ٻ���	fڥK�)�,5sQ�O��qF̎mRlqbXH��C�0�ZC�~i4?��f�uV�BϙE�	��}JQ�`��� �����hPz�����%F!��=F�B;���Z+-�{!��G��HN���f)�,�j�G�Ύ�GST��T��˺:g������p��h{!' {��ձF^�C�3}e:X���zo�[Il.��P���+�J_C�x]�Ϩ�)#����}>��گ{XT��`o�B��:.���zY���E�D�X��QhJ�X~��b����'�dv�veM��h�� ��=-�\ �����:����Ջ��2тD��>�o�8�,V�l��V �[���X"|ZS�.	{Ra ���b��w̯FK����E�(����^fP!�G>�Y�T�)���c��^kҢ��_(��P����,ρF� ��B���/C
ա�!4��� m\a��jt[�q����׻G�	�5��f�N�p�rR=��P�˧^I�/��>���N�������a*�ܰ��Bx$i�%Hff�M"�Z@lN%!K���yC�َR���^��"A���z6�W�n6ȜU!O���zl&X�Fp$�nj�p0m��l${t�x +���C�\iz�����6�Uڿ�6���%]���X,cc`Pz'/�:.���jَd��z�X���i=\�8(:-z�`�����Qv���ľ�K_�3?�b��8��x��xe ���gr�_��o��~�NO�oC��[S���b�~��φ*�6�ׄ�dKd<�
�\X�0r�����#ZMW�5��F�E��3�`bKء�|��6;�j�=j���ʙ�RR;�4��������t��iD�r��I�J횮Y�4 eX�7��H�s-9�%u�v%[3�g�~���\������F9$�ա,�.e��G�P`�N��G��um����vP�4�������P	Z�B�F7�D���!���"0��Cg2+��sl�tc]�C�
֜V�v����BX{@��
���K0U�:~}C-h��r;��t��R���řn�@_-�X 4@�Js�{�17P=th_ԩ�(��}�۰�]-N_L���)>��;ӿ�W?����ȭ7��'�����g���c����n�Mb���W����~�sk���H�0�Jc�!��/�x�޷���.�)�R��^ENjQN|D�έ֪�?����	9������/�ZtK�Ʊ�nN�}�{�3�>#��B|�=��r	f]��Wl^=�x.��.��S���j0"�`�X��å�CU�yA�ې0VB��ѯ�ބ�O� ���8b<�oT�R�w��DH���5�,��Y!קIbM�dW~�:|D=�&�?�ph�����ds�p��t{b�t�>��e�����C�.��N���-1���ZP�[���ҽ�1@��3��W�L�%��q{���z�"�I�ް��E-"���6I��\e��	�	���K�>ܣ���wަ>{W�yղSA��=jƫg��6/��0I'��
6�)u>K�}��ҹ��������^���4�T�u�g6�޺Fo3��Z�!�\E���6( ��:�ڠN]i�".���F����x�}�� h��(�ֻw����Ϙ�@���(�3(����;1eCF@�d�@�*��ЎJ(4s��������:�g�P���pگ]�ჇҔ� ��A|K3O0#Y����kYRk*a�tb���*�J(��E��ǟ4a�FH]F�����RD�4��n��M]�95����S��L�K)�aѯJ4���]�6x����Wt�,J�k_���}��Tm*%�n�t)�4 �=	u�I��룏�P�8� |��\����B� x�~&pJr��V��ϝ9�{YO���S�6i�;륅(r������΁�\���=�r�83eI�αp�##��������P!�5e��f��8T��fB�a�=.� {l��:sE�PHK�������O�
ǜ>uQz��t)��Z�VbU��ȳg��s��O�����l��?���;�Eao��&eK�N�
=-̥�g.lq�Wԏ�:�11M�.N��Z]S8S��Bt��9b��q��iR��Qm?4�hR�o��؈�P��9��4�=�"�S����H0��i�M
\�m(��*��²6�Y!�%$yYU�����^	ꕄ �2/'���z/}9ds�շ��	9�t�U�L9���m��/�=Q�0V�b=[ڌ�h�VUoHa�>��}�d��ҸB�=�I��C#b�$���;���	ٗ.MO�g$=���\�/ϧ�E �4z�>����~���vl�\b ���1�e�:֣^�l��kda기pu�n-�8�<��A������!{Ϩ��d:02�f4ޫ�
e�l°��t�Z(�Zm"/`��N�l�;����E��d���� g 5�z�a���5��[E��6/�z�>?�\D��[��� ���7,��Ǘ���r���bވP:���p���rwx��h��Q��#.�0b�F-vBQz��lsUU�U_�S���u"��-�K_u�A/�dU�_�@C�gT���B�w�P��޻����f�M���-�d']�4m�r��-�v
΍�+�t����2��I�:��`2x��㢯SM;�&Y`�nX���K�d^�t���wɡ8Ӱ��nBB���{C�u��]w�)0�ߡ��.�/�2�A�Q:�~L�k����8 ���[^ZM���:m�nxV����r��K��F�J'r�a"�����	�
�d��3ϼ�z�Ś��MKk3>��@�m�S�e���h����h$�}�b����h��:�S���M_��Uꢎ��f9�G%Խ��;��
ƅs� =v,-�Yx�;НJ?�o~A�ߢA]��]~ŀuB�=��p����ӓ�=i������L���#�>m}՘��q�(�p�4#����cj9|p��Ƣp�2�>��OHܮ�Ld+"���#5{fTaN��������/��
s�.�|��~0���gĨ��kr9]�f�P�=#�R>e��!E��;Op� �7h�ک{�O]]ivA���ae]Q��܅�tN)���Ǐ
�H#4��ZLoem1oǾ��t��^����(=����E9�p�knf���H����`��O��X@� �p�0k�#*k1��Ź�E�a�-��+��vҾã
U��[WAL�^"ʔ,����cK�c���H�g��/h�#�G�<7��Ph�������@��A��OD�K������0��D�^ �na��:���֠��1�5r�*���ޢ���&�6���������#�{%tJC�H�<�Z	������D�ȶ�r�4C�E�#�lT�Hk���=K�k�ֹh�����r��p壿�,P@�F<@�gAU�d��Bp_Ʊ_��ˡ��;�, �d]�f��Iņ�q�j�FqCv�0A�/H�7
�,k�S��_�?�wT���	C*����D�������Ϲ�z���W���Tz�v�6~`���4�����3j��k��t�X��'o9�:6{���%-����s�������EU�~��e1H7Yw�͏�8�p�L��{:�"�,�02�����4���~����s���R�ȣ��tn�ً>�1tQ@��^vcО��t,]����M���߸�w�r�O<��Ğ#i�7|cz��g�g?�i�3�^y�q�#��t��K�������5��ܼx�T�]ɬ0�=#\��yF�����B@�鲪2�t�tD�L�������ω�9cVbJ�Y��G��/�w:�!�c��^��s/������t��=�2�����f���y��xN��}D��ų���}Ea�i�/�A����R�d��������О��r�Mi����w�!1�z���B�U�>���d�x洳�p����E��MX\�C=؃�n�%�& H��9�6����^v��;n�-=��/:����':�%�)���L�n���˳��|N��a�����/�1O�
����3k����f�&^��"�C�����l$H�Ǟ�<��Э�{�=i���mب�)wl�pZ�|:���K��t%M(kk|r��g�{�!��=궮�K�#���i�BGp����_5�Tn`c����^���A=?bFHP���͇��ҵ��ɢ.fߖ�[1/��"/�~A��A�N�鬧[�H�|����
��.�
�c_���
dV!@�"���PԪ� yV��1�.����iI�NՉ�;��Wl��7����~��P���0�a_O���^��o~2���s*Cp ��_��tEl�O��_�5ϊ�����5�E�{�	��b��l�h� �p]n�C=0�I#���%� ��>;�^1�N���3��V���md��n`���S�Tw�U;34���5/��
��G��i���5?�o��'S�|u= b��b�9K�
�� !�"���ҀH,�t
$�@���-���E��&h$�j
�I��"6��wh��u(Ty^��KD[v���oI�	� ��$<ݯŐ��+�O�a��{q^�刾�;����R<N��u�����=��x�&�b�Ω�����E�>,�1�rp���M��=�,��
q�X�3�+xS���<:��?�ԓi��@���ǟ��q�^ph뀴)�NZru1$'t��% a�}��z<--	<������$��F���*�'i��Y�.�M�4&�O�u�E"�[��_T��lE��K�EM��7J_��w� J}^���M��)ܢ�0N	��ē\�	� M��(d��4�N9��Ys������{���B}���뜯�������ޔ���ߓ����#E/=�����KgӃ�zH�t:=��z�	��,���|L�����Oֶh���?>6��҂f��#��^z�Lz�����{�I�&) Im@L�зʾ�� w]�gK"�=���8}����:A\oKs��ԁ�'����Fk���M�y�"�*6���oV�W�ןx�	����u�l��E���z�g��5V��ٯy�{ҷ��o���!fQ��=w�cG�X�{I`��[�������Yb��@�P�r�T�Am�W�bH�H�t��+�/
|_����y��&ѵ X������{U�u��%e�Ix|e;�����ྃ���~�����z Ι�jl+P��x(�T�|QdZ����X� 6(�9��Ԁ6{Լ������d�� ��l)L!�:J�k�k��Z�s+�,V@cq]�IkG��{S���7L�����A��][���7���tif%�z�X��_������MiN�8�7���̃>�G.'K���zk")��^]fCKZw����%�ޛ�'�笣s�X���G�/g�z�|����x��@���<����?sq���к}N��0�X� ��`gۭ�����X���k����
Դ��J���u��3 +�[2,���X,*� {)6C �-X �C�'�'W��J��)����	�
�����f�mA(uSD�;kI��H�GT�b� �!`�*�Ǌ�-�0 X��[p�O�$�J��q�|�^�/��iPo���d����Pz3�\!��܀վJs����B#B��S�-�T�L97�|��
���Թ��[n5�N�����51���̬��ȴ�q�Ȱ8�U7s�"�%SL��$ȥ��Rck�g [��sCL�\^Ĥ5�	i��&��p:�>��1�'�h���U��qF�����N�O��.�� RJ@��t~�{�������(���'u]׃͇�A���$1�£�O�M8�= M�!l
�a@
��pP��4X�;�R E�h��~��#bY:�A&G��hs��ü��d	*�$�̈́X,� ���y[TH���Ɗs2g��% 
�}2oI�� ��ӽ�48�h&.!3�}L�1�E���Ze6�c�Ӣ������ �5 ]ծ�ܫY(��W���*��XX�1'��r����W0S
�!���(�,�h�0����#-�΂ަ�cQO�63���h�*։g�J�$,�=��Ç�:;�)�Af�������~�5)��6�������F��-x.�A���(�U��֔	�-��.��>e�W=�K
�]R�փ�'�50�����pz��l;v{ZQ�vM=�ԯ�W �=�JenlS�T�K�7n	�4:��LN��|HSE&b��6S��T�-(�"B�h�A�.�G�\��l���~����w��W߼��/Y`�/�"-P��V=JJ��nzU
�I������5�X$���N�H�]'���!� j���G��q��Wquj��?ґ������ήyJU{7��j(KpP�Z8K�}�C�IB��]�WBM�	@�{Se��:r�z��'c����h9�ye��j�cG:�P���j�Cs���E�Ľ��㡗�8�4m�USC����*�=t=� 5 (�;]�G��ͅs��TwF �].Α1bf��d��%��>�R9$����*��3���X-�
sىj���^`by�,����.07����G�u]8+z]�k��߇4M����5��P�5��@���&��Vz2�g����d���q)�&mz @aCYt��~9:@��3���2���bAp|� hB�3/�
��>����Y�V4�Ԉ!(D�B�W4PfJ䬸���H�<*�ɹ&'��"��ӂ�H��r����x�{���\fI���!���U/�<'�,'�y��]��͙�*HO��
�ҏJ8Y�9�{�-�<[��.Q6s����+�1"��Rr�l�"��%���w!�F #6K�_�a5�j��u�;����=D]�R󆐧�kc�,�HB��ss邴L�c��X
⹠�<E�E�Q�s\�)�rN���Đr�%�N@+E4؉��g�j�T�����E��zT!_����/���3x�-7y�_��r2bn/=ۢ�a3�ߜH�x�8���$s�RS�uv��w�s�ΦǵY |`J"k={�A1����0X=�=H��"�Z��� 5�Q�Blܧ~i�-������³���uI��ģt��d36'nz���d�u�=��(�s"�$E��u��%���o��nh����5�Ru=��SHVC�u�q�Y��P;�b�z���\�z=��n����k��:vCi0G�u�U,��s5�pL,Ξ�b<7;�n��f�E��iр��'�o��(��B[
���84�����/j� ���^br"B#cM	;�U�[b �  3N[6�D������j���M�N��jĹ&N������u�5 �Zd��ڽnlj��v�8V���b���%�?(x�Seg�u�z<UW�~��j�p~*2�^����k��rVїL�t��`g��Dqj�Ú����s��C������%q��(x^�*o*M��
�/ؤ7��)�77��@�_!A��4d�K�ӗ�h2���;�
z��jΰ.�۬a��6�+T6n�gB>���:2�)2�65\��N�*I/8.��QR!�|d��~p�0^+�WUÈZ38������cӓO|1���,�	]�4�#zb�Rd�E��q8kw���n@�ٶ��r��|�A��amqO���唙� B 5�{�5�b��I@��۹��k��3�g������و\��nXlд�ܑ5$[�9�֘qm�AF&�}U�Y�ߙ0Y'�k��V���3�ƥ�5��c���y���^_08�����F�>��%���c� �\7��;��.�#��( )J7Q��f�.������H���<?��ۯЩ2��i�;�7휺���J������Q��6�k�Ц������w?���z�K�2�6kß�=H�H�Ɩ�	�S8K6��P+�_iB8�En��Nھ�>�mK��7�I�!�Q>����#�]�@(@��=HdAٵ���J
;���/����z- ��D�e͐�	�U'Q��SL��ڑi7��L2���[>$'ؗ�y�Q��A��X�q �ä́�`Q\��d���珤WG5ޖ�a���������$`ҙZ��DNH[�B��V�Q̉B���a^�Z2cƂ���s����%�:}�;yt( *v�,�d��&{x���C	9B(-�2�U�F��>id�h��u�}��1' �� �Ь*d�]1eq�>�#��ġ�f�a�wT���'�	$��qЄW`��,���Z�G���7���ȱ	�^��ΰ5��`\�b��Þ,�A c��sƑ!� B�(s������CA�fg� �)I�
�ܙBUצ��D��=��l�������� e|希@����A��6�bh�{EY�̗��G�&�K�R�>v�(2n�έc �"+}Γ0�YR���ӿC��z:�(vP���ؒl  S����y`��f`Ђ�3;S=�9k���w�A0��ha�x~�!<�k�S�٦�X��J��mA�����u�6��L4 �eF�7���y݇�m
T���f�yX!69�dZ�w����?�ĵҎ�1䙀�@�M������6�>��������#?��Nec>��S����騴Y���`�$��iG$`��y��jp��Vm���WS=��{%�oJ�7�.�xg׺Z�4������1؀RQ������d�$����҉ae�a���7H���x���?tCc���ʊic磇hQ'�r(��H�%&O��x�Bȷ#�u�+3>�l^\�7�&s�����7��W�>9���w3ͯ��X�̈́��[�ܜ�������`Q� -���E��y3+��,�T��  p�cڱ���n�q���08ZO.�c�G,vktt�U�-��s�\�8ֲ�3�np����b�~��m�3�d{];� c��"���'c
_紨�j�A�;X�i�1qr:|o�O_�<�n�N���	sPtܫ[R躩��#ॶ��q�f� v�d�P�'�;y*�g
j Y��a�4+�Ыv�W�/�X �F��?)��+*�R���+'��������x�2�F�궉5g0R�S�0���/�̎R�N�ת�UP}0y����̬����U�!��9�j �K	[��+V�-j4�C��9���#����w '�^�!�M��q�{�h�mL���"�\���bg~�+�]tXp߯q> �μ��y��īR}��a��* �"�����5�r|7�����j	�2 �*�� d�L]*2�(�9�{��WWdI-W�{L�o�0�:6v�=���]��N��p2��Q����n�c@u9���]~�=�=�닁�d�	�ӭ�R�{.3/XS��X�U�h�O�&N�?��:#P��c�Z#�*��ܓ���V��ꏤ�nR�Z�^����������ߦ����tǝ7�����?}����G?�x���KE8�K7�h"�������9�Q��VsK�dӅ	�!��V�pA76b
�G����	$@��+�iS�±cǵ��*��x��M����3�^㕙�b^/t�+�8�6V�4p�m ���jw^���+��c�#vY=���P��agG؁c�T>Ο1+�F�솾_�BgQ"�%��?��MJ8�4#*��3���tt�'�=l�Q7��iA�,B�葚�G�Z�?����Q�/�!���\�J\K]L��������/�+Ph�B�	¢>! ��o��@��GE��ﷃ4��=�^P�'H���6��K�$v�f��w�jnݑ��� �S��\4��e�_,0�}#�� T?!0$��rxF��,�N�x�8Yvv�hR(9 ͔� ���$���,�Q\]�;h�0!(������"�=�e��0ЉƵnJ* [��D��J��s�� Pv��JC���*�n�j{Q9F(jOMN��q��z�|�"d@+�\\�6���95{W]3����A �h�g#�	q�Ց-�h��]�K`�hx*�K���ߖ�Դ~�V*� ��|g��+��QX��#�+𰪐@��I���_�5,篪�E��xƢ��������S��%�ı���9L]��-�mk^Q7,6��B(���(�#(��ϛ�̦�d� ��,n��4�k�1��CL}�=w�.�*z���1Ӝ��ZWVY?���--�)�S5��Lz�R�隵�.�|6�\:�nW�����?��u�Bjz��~,uJ5e�R��Ǜ�6��P�V��c���ּ����zMO�����n`l���ŮhH���[S[�!	�P�����E���z��k]J���g���Z�͋�w�U/���$�Ź��+��� ��+fح�||��F��g?����A��x�t�
H�����������u���ɱ�@�� 
���P�&��#�w�-��:���v�,�#����ET�p0-���x���]��+��A���z�+'S�;N��@�G��7������ٹh�\u;u��@}��)�������8 �1˃�z��~�M��N��2��Զ3mZ�XlQ�~�����A�
Y�*V��XTڥҰ�V�ɚA�c��]�X� Ж�{t3V�	���o�Oq /�J4��热a�Xo�{��Cv��¯u(g����fe;��`Ć��p��ꡕ�>�$����ju��^ )Y[��ҍ��U�ul;4H+4Q���|�!�Lc��ap͜ �	���������!?�=�3b��J� ��Y�=, ҂�zc�D-��
���Ǣ7�5��f"օ`� ��(�K�M7f��q�~���C����Y��<0��c"��7@�P�x1�
�m�S����W��k��䚂��S�j�bv5� �lx�n�!|�W���	T�q�/M����Z����	������2��z-�l�����c�k����CN���������/�L��o�]��u	��u�G=(h�K���"@�7�?�&]����<�dW�9�~ۊY��J�@A78�0�0r�������i���.,X,t���Z�a�|���ko�៵H�]�N0Cw`�������^	v��r�,�>�#�G�
����y�s*�����*�\M�k�A�׊���y���-�=/�i���H��=! I]Ǧx\�?��ԎI�w�R}�H�IKa40�:��]@�ԘZH��n>3`>2�B 	c;B�#Q��O�\*�G �:Cs'kl������gsp�B �
�Q��{�SޡFgm�h�ն�v�| '����3���}�Ҷّ�N��q���A9<Q1����_.�� ��k����>��b�pr�8i�� ��{:��񘹪X9dj� b�]dvˬA ��u-���GpK�,�������� %w��V�����ED�ss������O����~��p�\E��z��� ���sP1u�^��E�Г��A��9��\Va�G��?[��쮬!�Uq(v�z$2�"�	&�KZ�(y�&�Nr+v�Z�R:�8��(�����T]�5���h�|�+���y��_0D=fNSd{�06}�{%2�h��<>K���U�L��<����>���я}ʡ?qQb�g��魴Gw�T������ J��-F�v�*!�������O�gU��&���M��GT?죿�;��q���߭�PF�J�+s1�ɘ �h�<|M������x���me��nd���(4���ŋ�2�!�ƙ~ܴ8�v��A�������노�P�{ ��ڭ�Ʊ����N>����Ԏ�ÅAT������@����A(���S�����<D<�f��Wny7�Y��%�G��G���S���ZVZaG�%�oD���6X�lĪ���R��cf�q�;p�P��� ��[��"؃{qxR��wQ���M��C��w7�Y�>e�Iu��"�ܣ���Z�T�!�?����^�Vs֢�Nٙ16��|���<&U���T̀5` ��sTg'����a��Y�| 33 X�n���  ��z�TL�� ������!�Xv��(^HM_�O�
���J�gF�V�Tw�ze��	��� i�zs�߮��_�q�X<��N��
'�ōT��ܩ<O�;��d��
�
�G�*�/�\��/!t�W�' ��F!�T�*_`{��{蘢�+�J�(��1~�z��y>�t�O�; +%�9u��J�3Ĝ @Y=��-���~4h����۠���J�8�z@/�&��z�G��WNk�@�OT�����+�!�z�;�zS��U�?�$��
MN�ێ�ǀj)��gYa�Q��P������>����[|�*M�j�0�ޠ��[���0k�ϸW����6�Z@��]�<R'�X$a%H&D�߰��@8���ӗ��uA�70�ޟuA�y�^0���9B]��Z�w8����_��_C�gRi�CC���=�]��� �%�Cw�����iŅ�$�`�Wy�_�8�� ��.����E2ĴСu��:�ߡ�!�-����L��n!D���J����Z��S�A�����Y��G�T��E�AF 	E�2�tH
A0�S�T�=^L+����b ��lv�E��札�?��Q�$�+�fj��)�r:_ճnU>�!�D80�f�{��v��X��g��X� �h;�*܆�B� �@��b��k-�BQ�i�b��D����C�D��vE�b��e�+0��ư 3%iM������"C��P�u`� ���eJ4�\�.T04�˜EU���r��.���2���s�9�s��=8�����B۳��V�b=e{�tm%��m��.��Z�e`�Ƈ����&�/�b{i��Fu�j�dMZ:zg��s���1�L ���5ޤnU�N��<�z0 k��;����NY];��@g�l�P�]���$�� ���Kz��Ҡ �Z�l	,�m8:qo��{D�ɶ��k����B�ϧ�S5x���ծi����U�W;�餸·����Q�����̛�py^�y��o��/]���/_�( �؋�!2���B�]$R42��EeYB��y�*������^��}���b$�~��, }���xy� �+����G�%a"�s�^�ݳ�=�N�<�+�ʎ�k�I�C`_�E�(.����G�+R��y�v��u��B֖�MD��OX�z��5g��������&v���8\�0C*��r/5] �!���6-�Գa�cLO,Bh�q���w�Z����=��� �/�Ѱ?/��_ΒB��3����1��rbLpN�3��	ge���˘`[�2��?-��d���F��x�tXW�<�Z)������� ���p�<
��$������b���b-64Nd�p��A8ƃu3kU7�Jg�)L�k���N�ah�jNȆ��\ȦZ�c����+c�0��	�� �^�����<���_Fx2XK^����'ol�� ���*8����d�t)Y�_� һ�`P=���`�u���pb��K<`���W��+�Ɵ뭴B�����D8�Ў�an� }M���e<�ޔ��1Q��W��-��ੲ��"��V�2
*R� �=��	���8���e�9w�!�qe��U���ǞH��P�cbxb|(��-����H/����S���S/��o>���C_������>�ZHL��6�VT�r�[����~G��U6!Ɨ�[��D��jm�`�aH��Q�!�X�</�_�m[��[����i�� VO��m�, �Sv���wd����j��m8vw���/;�|��s��p���X���Ñc�X��ي)�n�b�u�e�}^8��[c�(!���R�O���ϸ�Zv�A���Rz,��w��L�7��y�ov"�ʐ5�� �0�=@���~pB��PΪWY0�I���3�Y0�/�uX�96�C��q�슲m��W��h�����0��E��"/��ٮ��������[#�6��m��Y
E�"�j�E8�T�(�3�xy̮MR'���}.��Dx�q1;���yFc[�	Pv�!���c l�K�ܰ��b�]���w������}��	��}f����a/��P�X�����7�RM-;6�X8)D�����z��쒾���ܬj1e�n�f8�e������+>����󳗻��>��: �V�h�0�+Д7j�� &���&Ѻ�HK��?�"�0����{� ��� ,��9�ˡ�T֨ut*���me�u�!�ҭ���[���M �b۹:{<[�R���������Y�Ϛ��;�����U*����~�JSx�Jh�=c%��ܯ�aSz^�g{�e�5������Hz��ϥ�O~:}�7|M�����a���H{հ��3�%��]�.��R!͖�9,&p}��:��fgws"�Ҟ�Ǒ��H�`m8J޾�B��sX��ʱ@A70�b����Dvj�Z����a�-��wC$��\�rm����1�	�8FZq ��^t	����T?
����?���~B�wv�~���8ip�[�H���8q(htU$�2��}�Z�n��v#(��"Ev��v��P����C ��DQ�������0A�; �$=s��$�uW @�6,�؂�3EϢ��rc����^��1��L��rj�r/&>��w��ϬL���AH����$C�0����c�do� ��Z5Մ��Ɍ
JUx�c�6�� ���@P��F�}��0�ò�uS���!b  DYU�dν���`#B�l�g� %g��T��|UP�خWc�]hQ���d���ۊX�E�b�6���w8Xq��ae���E,����2��L!Ć�'Bd�x�0hy���Q<S{fs�У��`�w 
~2�J�Y`@ ��I�7X&lN8��"��r�ޡ8��f��ɫ����3�A�k2Us�S�����}���� ]�@��F���흡��`5�2��a���\���w9����L����o���BXqe���>�5+�k�I816����>�9��:Y{�y�"���|.�-�N�S�ĥt����g��;�D�f��?���o������f␒��*G/ϜK��b���F�[�'�֮\H�c{t�z��.�a��"k��(�bW���W%z�yh�vTF*_�b-P@��ŏ<�dh J�	*'��v�*Ȉ����ݰ׫v����Z Y8��)_c	�q\,v��+����q|���� T��w�����[hГi3(oiX�F�����p}�(�F�`��:)8�\Z�EH�+�O�Km�N�#3X(�ƚ[.�7�X2L �K�$9/@����r�1�i���p9��a�pX��ݱh�� ��w���"��n ���g���}1_BZ%
*������b_Z�-��:��C�N���T@�V�?�F�v6�Af��5�}p�v�w9ę���T�-�����z����P������s��c��k�=�dܶ�4���O�;�!y��kO�ϟ�kf^��:6a�<g�O֥�����G����,����JDϥ~O�c���}سhIr���PT1�c]��d���|��+��L���W���b�}����^��m���@�ȿ�� �s�H" D��</�^�r9P��cG��)�R�'��&�k�Јjw��r����<���ȁ��?�G�?���N3ϥ��qO�'�׿M�<���J��a��?�W�w}�itl ��?�'����ӿ��O�ob'�y�0 쫠S���bp�h	�fr�Z#:{<vz��T������`{�(�D�t�~��ơ琉����k��ݹ�ﳳΟ�#m[���*��j��gX��
��� ��r�.�c�]���w����e;ӌt�l�VxD����P�:BN���v3�!>^��d���Ǜ�V�� �;��8qt2���؟�+ʎfTUfI��E����p�.������l����B}|6���x;�g&%t!�_ΔȎ#�K�4ؖ\K��f%8��#��]����jg�vME��]xv��:wY�G��+g���h�dp��(�;��2 �Ƥ�g�\�C���w��/�J�l�>��=gJ�����אs{j?���y��8��j��5@�F���z�����"���=,WU@�kʡ8�*Ӕ���ڀT�������̸0N��lg��}�5__�e{g`���������E;j�����Ξ�s��l���pc�?2��!�&������_�m|:�o��� e@���N
$I�S�V&m� g�ZS�U�`e�R���iY�g�sګ�?��%�ӟ�����1Z�<t�	�W�Fu�T���w�'��o<�Z�
wB�-��-��Ԑ�󘯊�Lj7�v��IL`�T^o't��J{vA<M�2��Ȉ��o2{�z:���Ũ}Qs���][��]�S9*��8F6���'��Ŕ��"w�vh!X��c�A�+07$�Uj{%.�h������o��̠�㤚v���q,.��G����ݮ#*\��z���i!��P��δ�W�q�bprd��{r�C���uBUZyδ���`�||��Z�ɋ5�t��l�v��N���%������w����PSe;Gb��[W����k	&��fdG�=��U�ZT�_;��E,�|F0*`G�q�]�3���<U�I�f���������Y>O�_��8�R�#! DnF�_�u4g28�X�@(_K���}�2@����S��X��A���b�2C����Ӟ�9ڵ�ϣ��lH-^yN_Ϩ������Ή9a�G���r+�/�|�0��$V���σY����v��k�6kg��!���:!d�M%.P��[k˅��s�=�z�^_�������g{C�������:�����ӿ�qi���&������'T}],r�v������Ks��JX=�������C��2�$��5����C5h�:)��Z�X*��<n�ύ俜�\��ֶ@A72~A�����9[&��*QB8a��^h�䅟�U%��`�'c&S�m`(�C;�l�Cw�M��~[do4�k�9��z��%RdQ��d&�_�bݍ�F��c#lT�Z10?�?�^~���o��2�,/n�}�rF�C3�"���]�v�R9;Z�M�?���I�Z��G�\��3���(h1(B٠��vod�j�Ɓ���z�B�%��0L�E��#L��:��x��y��k9~�w�\��Z&���Aq���ö{p�w2kD�̙j�Ai�σо=\z�p��<�# �����^�Η�v������D/�-�>\{�厪0bv��[(_��<��9���<��͈9H��k)��X��t���ܱ����g(�_���/^��l��L�#D������u�^ZZh.�Bׄ��Y�L?>ü�=��B�و��q���<����t2E����'5����T���ֈ��u\}����\��x3��{��
���q��3�m ���y��I�;����F6�j�#Y�Z�\1Zz.jt����>Uվ�������m��Tk�.��첢=-%V4	�S�[H������2�������FLY�U�jC6��Bz�����+�o@��c��m5\��I|�u�[��~t��ŤK����k�p��GJB� (ov���W�
����Â
�o�U�Z�^��B�Pe�x�Ks���f��n*�S�+;$��m�bU$�XY�I�]�r��S�ISo�MB	I�0� �Z J�8e�ә��
0�:��}����N�N�v�`n�L-�Ut<"�q= �@tnc�����Z�Wɤ�D��T �k�K�CF|Ζ>5ObQgA��C�s0]�fL��*������<q�0-v8h��69��w���|�<��� ��?�Ϻ��w�9�9W��1��2���l��=J�'�M��EA� f�c�(�r�^�P�'Ӎ+�˅�48���C��*�s�,�\1��%���Y���=�Q���{?�a��!� �U�r����~�#��Ρ�0�ưC��{f&�~)��s�a����i��$����ɽ����0!p^��z��g���x��hZT�΃�79y��ƢP�։f�yn���������-gp�pf�8e�9�Ky����P�'�J,\o7�ٶ�p��z6���*�]�-7I�Xi)�>��j��GL<���QC\���^HT8q�ѩ�óʜ��3�uakD�qT}�Ⱥ՚5��GBt�Ue�=�S�(����t�5�e뮫���O��ށ�jk���w8�O�(=���ɖS�j&��Y�[%$���+���n`�]�ǆ�k�����(�H�|�6�v��� '�ȖKl�5�E'�>߂c�,����V������E�`/��m;�H9��7�ќi��E�ؙ��,k�1�	zE�Z���@h���Z�����,�)�NV��q�
}��#b^Rh�3�H	A�.�3�T
�vyv�0/f�9pO�~P�BdS�ɺ��j�}�
��8�e ̡4X��D���9;��1�L�흮�ag�C��}�踕���5�Y�p8��r�j.U�7U���^P�Y��"2Aa�.�@s�Kۡb��r�9���a�k�s���qf�<�"�ʫ}��Gȶ���|��jKgǜ�'��u�T���sw���9��������'�S\��!�LŜsH���Ffo�D�&나��ޓ0D��������2�k�z�.��'<����&F�!�x|���U�W�Wf�4��a1��W����g��EMK��rTѮ�:�Cy|�����ꁹ'�Γ���S�и��y�WZ�.�p�4D���IG��sZhc9����t�-��w���H���w&z�҈��h[@gG5�:`�7�錊*>��K�"�]N�lߧ�iSi�0b�Cc�1h�S�=S�il�xz������ϦgN�u�X�޳���T5��̺��(���.�{k[���7a��QTl����Z֑uBժ�~j����WC�k�}9���p�_z��Uq��S��^G�{�� bfF��A�!����bC|H;��z@�j�T�e�"x��H�%����Uub�wC��)�hc�ʵ ����)��������q/tg!5��������n��Z��* H؂]7bk������>�� Qt���\s�F�q����O����-[��i9sث,"��q�륪a�Չl1��}~�C���4v.�K�&�F�0'��Y�g��cG�8�qW��A��r&`u|�o.֗{da�-�6�"/�@�C��p�赢�|�+��'�z����}�2�j���Ɏ�g�7 �����p�k���R�Y�� 6!�e*�ﶁc��
��T�����v=� GNq���s��0&��k 6�箻����64�７1�S\=��)�8߻Ǩ2fhŘ/h�\�gו��"�.������g�eXf)��.�s�{Ό_imx������	��4��>3Fn��zAhv�ldd�R����{��w��Kcb~'�G�g>�4��8��ݷ�P��B��?���@��;n��J�h�߫jLs����ڊ�"��-b����)qف�o=��<pO�V���z��ОT�<��*F�n��Q�^I��Q��L���җ;���ߺ( �Ʈ*W�nC���\U�#�A��pp��_�I�]���>�ŧ�3�_z������9�+رR?d@�b�z'Nx,RU:&��Ml��X�@�]g��=��Mqo8�\���a(m�o��֕��w�(`Ȃ�N�0:W��"o�&G�K΢��PW(�E�ir�ܢ!gj�� ��\�k�εJy�ޓC/�/U�%۸��iw�v�m8�ރ�u�����3��]!�������{J��3��H[ �H��z|e0�GȩЕ�Y��,Jf0��FA��dQy��sD��1��= $1��C|��P���7�q�dV�}����Ο2
��$�2�k	�G"�n����:v~&rh�lY�2�[b�۪ @�_>��� �
=y|�^�N�2�`;x��O���z-���1���ܔ׹6�s���2��#h�V�l�2l�5�����٬ |���Ҟe�{ܪ��̲I{)�6k62��*�)*�,H�M��N��4�d�	eq�x�c#B��U���J��������������[��c�	ZO����l����c�~���4�sZ�۫�Ѭ}+�J�P��m����|z����<�zǦҠjK�=��(�ZE*�RFj�;���@�'��r�7:�����( �F�O���B�YO�cY@�v'V�W��|j��������}�K'r�{a9pZ�:i�.�� �P�MgW�R,��e��*�2�X0�㇓��[A��{v�xQ�)�B�+�Ąi���=����1S�uX�Va�c5w�X�V�u=���g̰T:��H�����0��]����sv�����dX<�:���F��s1��5r��U����_�{�ﱑa��6���3 �nt�4j�1!R�:,���u��s��Y'�Ӳ3����mƞ{��'9��E�@In3(əKo��ɶk�d�o2X��Dv�y12ۘá\C�c���� +�7�<�.g����A�k-��p��e������&&��Ŗe]U~�x��_<_�����E¼)�]/b\�}3v�;�v��J���%�N���y�SE�����}��h����)���WM�c�!���Ǽ���y: Kd�*³k�K�Ra�(w�7~�7�G�|z��j�XYW�c�;x츲��B�W��W���z	JX}uz.]�zE��H����耲�.��J��M������SuX5�:h����u�ֺ�O#{���7�ڕ����5�u��|m��"ݽ�8�v��7:����R( �F�+�UZ7"��A��c�nn���r !^�lMv濙bQ�V��d���vГ�z�nU��k�Ϡ�pJ(�Cג��P��Q�:@HN��*���k��YK���ѫbuz�e������ ZZU�C�C���Ř�1@:O���l�
��b�?��_�)��4��(�2m0m�����g�9��V%
#U��2�$P
��@�1��l�G�uL^��W�OֺXoD(���haQ1��i;3��З��~\��v-�ru�.1f�S��,ZdD(��{[,֎��l��Q���؄��qrϙ!�N,��tݙ�����t0�E�K�������dp�>gہ��\{fX��8Ute9�
�GO� ���=5�9R1{yNy>W��^��*t8١�����C�]f��v͂��3�����e�����+vK.�Y]���sߖ��+���D'�1DCG������wD��vf�k6���=�f*��5�#z~�Ħ�V��M)7�}������V2Ӫt`���0o�UC��)���3�H���=��`�V���Yg�޿_��GF�����)ė���H���P���� i�N?��G��.���f.+D��^c{�hyM�ohCﶦ�w��M}���3�����z^���K+�*�^O/]M��t�����J/]�����*2��Z��9!;2;k�}9�[���� �aN�5���o�X�5��� ���,��_,�uA
>X�W�|�ICT��w���0܂�n�z�1gMƓ9�}u;yb�ľ"L[N=R��.�܎@Y,��.ޘEW^P;����N��.40hk���ڷ$h��`�6��4�ۢ��@߀T�uD���Jݷ�:fcv[nha�q�d�H�����Pz'*튮��#z����7Ů�zk3hԩ���0�*���Ԕ+W/,/�!���+]�#���]�Ȣ�` �	
p��]{$�CE��*�X�~��B��{tMjsВ&�~R��DcXgV��z��"�2��l�a�3�3�<]3��z�U���U�� Ե`�B�0A=�n����XON)�#����[ti���!1.ن���Fֱ�@����=NլW>6,��� K��m�����X�e��я�{U#&o:ܚª�pfܲ3Bbͭ`W*��ff�����!\�V�0=λ����j:�k�ޖ�\�Z'�K�]���*��#�HQ���W�&l2�l&�,�Ě<3���	P8BH�gW6Y�Ƃ�����a��h}⢄�jγQ	p�}^��YD٢�����CG<�n��k!�ݛ�{�Ζ�86���ٳiAa*lb��6��N�s�Z�� ���OC��;�Ÿ���~!}�?(1�������[Jm_]ZI'�I��#��4���"-@�o�^�G�.S)�kLU�WӲR�;d�~��U�&�t�N��.i�&�>m+����t�i�؉4<�H=�;;�Щ%�m���j��64M_�������߿( ��F��j�"�ˡ����*ڛ�k�D�|i
����.9Ț/yw�����ô!~�.f�PJ�-�C�Y^"f �FD@�B���om���ڵ#���{Mяǎ6j�X�]�`bWkڞ���-C#ғ�G��r�ⅴ�^Qd���S;�ɀ(�y1%_�o�T��*�d�Z�oto�>�y׍#��[�NO_M�OO�Kt��f@,���
5�A��W��i7U9\�!�ٱ�rQ�и����-̾H�	p��.���dG����U�0��"k9�ʑr<7��f�SV�O��S�Ք�&FN�ά���Q��?YKE=ܜ=Vμ7?~\;�%i9f� az{w,v��7�������-s0��x�Y����"kX+^�|��)��}�Cfb�#�fM������;�
��53K��c��RT��[i��l���0�1cn�&��܎ۣ��}��F�sW ؙ��]0���A6+A��˕7��g�:\�bZ�d{J���o��oN��}�e* ��S�BsY�o����#���du;�������PGJ�%}sm�w����!B���g>�~��~L�X�;��-�++���]bnв� ��U]��ŋ�
�t�]w�!�η��ѣJ�2�h�+0pb̯^�I�
���t�7Ž���I �/�=[N��,�7{媎����oJLx�*fh+�6WӰ�*����Ӓ�ua^=��6Ԭ�G��Rw��N%�KȤ^���j��_�( �6H�G�	�uo�3��W��p$�<�ηS�E���T�8�����رq�0"��8j�IU�Tv����~��ZY�0�k4y�1�D�����p�Nd@�ܢ#}d�D��Z:�w��}�{M�gMC79��>���*�߶��u�Z7�f"B[����2 bAǙ�����Kit��n��Q�`Ɉ!,{�`��c��m�h��-����XiQ�r�]���p�r0R�11]��zk��?�i���Ύˎ�� Ӗ�qe9V�l+����`��М����9��q����}�;#�l��r�^�Wr�^9J�J���6�`�^�ۀ�'6�T`C�0&�	.���������w}�w�f.Qp3�$���x��y�����[;k?,Snw���7O��7�?���@����-k�r�0�١!�6�fi&�o`H����|�ؘ�ߎ�̡!9���]�zw�_��#�ߛ�������Ӯ+�&��0<W��|N�@a�{��y�	��ʛ��}��;p�������7]����d�Ǌ���/\�ܿ�[��Z�%^�银"@G6�#�<bM�7~�7��h���F��6Ŷ��ы�@E�]�1�7���@����<��X_z������ϷZu�s�lR�gGzƁt�������l35S���k�4���}�0S&Zss���#�z-���
����Ro,lD���� ������]`!p2���%��xs�+ǥE��ͺ(m�U^��3�P�:����'ӷc��p���Jt�'�� �����Q�P�����*������_U;��x�0A�D��13@q���bސCw:���[�
{ 3+� 9N��`�^N��|_z���ipX;X����	�  D���3�K�Twg�!��,�`uwm���[������p����O��?V��;����Ä�e��9),�x3*�ŎW;`6��a����lH�2��-�}��O���O|"=��fw4��w!ʪ��+S@�-�P���z5���$�sc�X�C7,&l���[^I�|�C��sߟ��m�e�t�^�K�.�^���Ei���xv�j�|�v�L�g*>*��� �(4CX	���ރӥ�p���59�V��|��Z����`�ٜ���PS�I��n���tp~�#j��mzF��[��*�6(M�$W� d�E��^���t |]\T���(�������.\Z�3����y �����?K��P�z����=�q���}�������[f��U�bC�u���[�w�T:~􀚪Ω% L:����sS�;b�-���v�jg�3@���
�i�6]��i��1b�R�C����s�!����O�m���"	z��"L�X��?)���Fmg���e�&( ���sx,ZZxs�=m�<���X�_ ���_Z���𲣮��)�8s.�~o�A�'4 $x�i1����t�}�Iԧ�⊳�ܺ0����u�2*}�'\�g�ӒRsYH��k�&}��|�ŨgN��uf�s��ώawW�P��a��w��E�ŕ��
[9�xo��ᵤ]h��[T}��j��#_��`P�KQ�:��[�ȶ𢻦ٮ��@C{K
��`����w����ZD�otIPuݙ��3ϺFM�N��0 ˵e�c���,h��xe�;��4r
�y���4�GB6�����O�9��^�v(���뤩˞.Pɼ�ޭ�i>l���}�]�/�~&��9�g
�����Р+L3';|�?���	q'+mJ�-� �}���+S���#�vɀ"_weF��Ie4gR����	��^I�o��t����ҬCG�����R9�����ML���8o���f�w�����;q�Ҵ�9c��c_L���Z��=����^ �J���m��	�X�j'Qu�LP�Q���V:
�nT�G ���s��F� A�U6��r������~��ނi�c<K04 �?�?��t�w�Y��B^u�J��K���+.����w>��i�Q������1�����Κ[[k�q!�F����W�]��ӽ�ݫPۢBi���Z¨�ز:�SChyI�[5^�R��rZi����v���ꍸ����i�ʹ��`G������6�@A70��o��;^���ڳ���k�������@�|c�^��^��W��y�� afK���%6[a��dĳ�8(T�D#�LiC�9���#��8d' "L��P�3�d}rT�m8kI.i���l��_x����w�ig�vf�lvh��?v���v��b{��bQw�����By�f��[o�9����w���?��:s�t��N=�}=�B���4��Q23���W�A.��5y�����,�n}���Jw�f�SO=���������-�����x�w�a7�Q�{"ٌ�Bt|m9D�ٛMi �4+�O'�˯�z����OX��cv���-G�� �f���B�U"V�-ɺ9A�+��)\�:�^�������ΨH�%�|~����������wλ�T�F���v�0f�=Ö��"ff�~ה�h�Wd]99A�0ٺ"�b�������x���?o��o����!�=}���������ܸ&���A�������Y���Z���a�?�����J����t��)����+�����HO�8��`�t� �&�@�wg<JϷ�Y/�\�~��Y�K�B!����N�^�2x�Գ�6�����Q����|������~o���|�����=�d��u�h�Lv�6<���(�}4�TK�Ad��]��Z�أM���\�j@!+͛˗.Z�`FC����-��r\ӈ ك>�гt��	����t{��J��Wl���}�/}ʎ�@�0�G������� Ͳ��?�cwUu�ӓs��f�����` Ex�
�$�$A	��������a209�ι�+����}v�3=��L��?�z�����>��{ιg����{7��L޲�o�6z�����p�?���ge����A����w�r�P�Ŗ]��r�{sq5��X�@po� ��c�GcPŤ��®ҡ� e�Z�>�b�2`������V���92@ۖ�\c���gE��ػ��U��H.�}j1���pQPv�ZV�n�x��y������c��򒗾�|�/?PN:�$-��eb�ds�w� �����iP���Ge��
������Զ�2�~q˽���QI���>o)�׭.�~��ʕ߻���������m`0��7>���?���n)��0�O�� �ņ��н��/�+amy�{��0����1~ի^��o�fRk�L���njdD�8����$�7�f_�%C��Epޣ�>�;�O|��C�Pٹ{Yѷ�<��*O�姗/}�?�"Qe�"jǟQ�Z�+�i�Z�iD���dL9b   �)�	l#��)a�Qrý�o����7��|�ӟ.�wn� �����Cҙ(�7ŵ<���܌$Өsdcj�`	�yWb�v2�;���c��s�5ה���_�˯�ܺ��=����xy9�Q甯~��:z���M���;٧|~���9_y����F��������]��� ���\nP����9��{��_'v�!EG�	L7`��)�x���"WW ����ϻ�ȕ�AkƆ�,R���}�|�ӟ�u��Fz�ﾠ<��Ow�����7�7e�r�0��D���Sc���zѧl�\�c����G<L����>�պ<~�[�^�֐pѹ�46���ͼ�����K����� �� }`|o���r�-7�1=�]j����A1��{U�LݲO����eU��H���vn)�z:Z��̝�7�y��̎�_�;�7�{�䁡Ѯ�ˇ%؞�Q�f�=oko�
��sV?3�9G�-]:%	�)X斞1�0���w���90H)L/k��ŶM�)E�Y�ҠiV��g�:N�d�8��uP�]_V	��	}�ލ��ض���.����ꁀk����	�%s^�{��u�гkqqH��N��Hj��EhQ�"����"�� -�]��yR���{`��q:Hn��kWy�w�o�;^�6n����@�>�z�a�)����_�0u@�1Io{��yQ��<X�_��xg�n�7�,߁�O��l���^w�,�\�벀��q���AC��7)eㆍ�������(�Ʋa���w���q�Y忾�������Y�%�'��,0g��yِ�����aCW't��܉��-�|�3��@ h��QY]^����a�;��������]u�gZ3sZ��l`�6퓼��5���6�ȵw���iW�x���'?Y>�5 Z�r���}�s�)g�,W�x����]�I�s�2����R�8#\�b�9���k�d�E5~fA�
�x?�)O)'�|�������s����r������=w�`՗�a#R��1�Q� ����O�>i��G�t�l�pls����B��G?Z����ҫ�9��򲗽��Y��ܦ�y��u��J��2A���P S&l���.��VKP�X�:>�3=�.��2��8���EP���-��|}���?���=��e��NLC�O�A��M�^}f�(�`�������:���7K/����/��^�yĜ����ny�����#�K.SD뀑��<9�)���a0u��H,{�'�sĦ-t���Z�tTEs�ca�����j^S,��DX%�L�����i��l����,��T��2�	X�j�-+�^zi�v���7/����S��KK˃�z�X�����o,]-�=m������ۚ������ͱ��M�M*tR"r��5���ԾwF�ш��P��wN F�;��թZcg�'iV��h�פ���r�c6����bKZ)4;�ci�d*��tV�lLl�>�ߴ����;{P}�P���5�����/}�.��9m�O=�ԫ�>�+�CM�O�� �0F|^c��P��{���;�{[$�������TM{��6<F_#�K�Az�F�(!��wP�n6��,�?�9q}.=��d}�Q�%�d�|��֮�B�{���Pn��E�*���b�0�0�$��A���ǜ��^_��W� |�_2��7������/g�u��$cs��+|<�m���*�n���
��ݥ@VÈ��}�{o�R%���N?�m8]�������=H�y�\ ��B�Y�@Ȼw� b�Ƅ�h��~���XM�U�N�K��q���x/��r�]���w�׼��e���2�������=�l:rS��5�h�骰��1}���_C����#�������� ����rĚM�w����W�W�9��[�̦��B���d���_A(�EEe���qM\n��	�(��E��42Z�bæ��S$�P�z��c�)���3�]��������UX�𕯲�Ρ����sA�O2��u��'P������%[c'훘+�͜���`�MoWoy����x�+���!O���;�0� etW^�=�9��w��R䍉�B����R��Ѳ}�v��?��﷼�-n��뿖e�׫4Ĕ��p	�O�*�n�p�gA�y�Щ�c�o4\qfv�ϸ����>H��s�����?��.�eT��]��qDs�R%���r���[��5��h�y% �V���4����l����vq$t$�����:�`��� �y��Kӽ��%���=9W�"͇k������H9B�չ�>�\s�5嚫�����	
��9X�%�����꯾�%e�e�ms��g'$�l���kmk�`M�RL�S�}�\��w��v��ܬƱ�t ���Ҝ�̜�g3��3���xN�����]�6s:fN� �&m���� ~��zf6�75����Nj=��'=��#6m�������}����_���0��O�WA�����4�zḿ������{�EŬp�n�mz���U�'��~�py�cD�G!�3J�7I�0��X8-R�y��6Q6��߹u[��p�)'I��;|��K��c��I�T ̤�\nZ�"��6U�W~ �R�u�7:��Moz�싾s�������򗿼l�$���3wև��7�\�<9ћ�w�t/,��;L�������_e@.��2kN8����w���r�)�[n1xs^��%8d�%�^�}#�<������#�wja�'랓j�;��)*m� F��IO~�ټ?}�[zv���ۿ+W_}MY�c��$C��z��  z/rN�d�</ݤЁ`����X�p��6Q^�◖���۠n��b`y����o�9���.J
�6�~�H�9	�i/��ߓl�e�&��dKg�FRu  !*�2�j0D�/zы��A�>=��o~.�k�xq>�~>�^.�&��ZTXs Dx6�,=n(��M7��{�� u��@�s�����?ݶZ�x�]�����Q_�:"��$ &z$\���G���Qn��A.B���.�`�φ�we��|�Ϲ01�_jX��g{k�2�9�b������?�s��t3[��J�2(`@j~�8�21;�l�]J�1w���r����+���kָ3��v�~�DKp3N��]e�`�p�"�_��֖Ve��͑
�Dݢ����u��?��;-&�r�U�/�vl-S�=*��?���x�1eǖ������\d��Hͷ��+��ڿoN�[D�4�uv��u�x_��5I{47�bE3A�<��rF��Ts*�ɵk����Ӥ��\��m�C}l��S�6# #��J7��A���o��U���9�E!��a}4�N=����O>�G�����M��}[�]uǌ�ϯEt���b��$R�i���@X�{|)��=�?tq�/&�����y��ު���3㢡��"��t�@����9+��E�J���&"�N��f��M�s�N�u4����B��%���+F�W�1;��2��A��-R�<8(��}v�K����b`q��U�Vڨ:^�җ�=����n���VLǰ��a�%uR��
��I��2(S�!l&[�������Z�I�v�j����K��h7.B،FÖ�+�q��V�)�b�������q)��(�1�hX��*_ Ӥ�\y��~����������f�?.P������UF�j(3p����M�V8���r�/�vW ~"j�E��v�1�KUy�촓N���V~�)?�]+n8�"���v��A��L���E�6��(q��\��]��=�E��Ι�X� �8յ�y����c0 ��8|p��)T�&���|�����=��]�Q�t��oZ��
�ݤ�C�D� �I��a���]�l��K�� �
���ҿ}�u� �,�Ò��}Fs�%�����W��k�q^��g>�:\��I~�(l).j�W!�i@��"e$N����=�صx�:�X��|�7��ՏU~ƅg�1Kw�-��O�y>��~����3�>\+F��c�ZX��o��\|��z�������[>���T����v���� �Ѯ'] �_����_�)%q"����g��eҰ��,k�u�c�*M��u��zB�����ȁ��n.����̌�<�]��jͪ=�㝽KF���)Bv���D����.���葇wfF �S@��j.��y����O��aN�O����j�Ӧ�jQ?�h l���6������S��K��i�jW�~�7B���u-�7u�c{����ƢYk���'�x�>�G�C>_A����Ԣb'��HZ���V�k�w��K;쵨�'l�yy�3�d�}�B_Y,��1��,..@FwZ6e!�H�ء�|� ���916�ZX���.�k���Yvn�M#����2
{��uJ�=H��=��`�5F�6�rqӈ_��|���[�������W;] z�$�|�+^)V���;���ZL34=��Gu�%=J�z�;^���Y��$��P2�#T=�"�9]E{���4>��L��駞Vv��N�pT�۬E���Q��ɇD?�ֱ��q�ӎ(��;Z�,�d���C��:��(Na�P�N )��s����/~�\w�JMp��ĥm�;�6� ���5+�8�>B�N�U�)�Q�"/�� y��Uv/<��s˳�9��7+�x�4'\����-ޠ��2D���u�"MIv��ġԎ
�t���pM�t���U9dd�	E9�.�j"�RL��0�-�H2��n�Zz�'sSOh�`	8/._�`�hDJ2/ �f�@̙�#�U>W�'�Ͽ͞�?\�������D�x�1��nW����=
�)U�9�Gf̘/5h 3fG�e \���ah�������@߀;���/������1�^_�� �+�J�ad��H��G�gua����U
@���ث�ӹ}t�۴� W��MG��Qcܛ&j�m�_yy�=�q���//;u7����/~�<���v����F$�)�x��6�M_̨� �{Cr[�M*��k_��ǋ��㞻�a[���w�܄�Q���t��^m�Vo(�.�:x�ƳM9�V�9;E9��^��ѳN:�?����(|�U?���" ����M݊xY�U�����?Z4O��m�{V{}$j\��q�G�9�$�����uz_O�^b�[�<�]�ڪ睷c�B��	��t����3N?}��������v���zFv���s&�� �0�}fl�yv�%U�>G�y!0v�'�C2<
cB�{�X�Bg�lR��o��g���qP"1��5! D(�X�v��e}�on�
	���U�hQY"��Gn�v�
�2d����d�D?��*C{����yO��3	�z�����S�l]���b�^E	�
�/���N퐹=���TbqB�D�!S�j+�vьLkGv���)c�F`��J�j	i�c�B���U��->�]e^�CTvC���
mN R�����R���qF�x5F�y���	'�\�ؼ���k"��KYF({��([�f٣�b�����Nډ
Q���ݸ�?�o�S?Kd;.W���$�,�BH)0�62:]� �}h��N\��1�2!��\;� �qjfL�$ˮR���Q_H��p�EA��aZLaP���M��'�~X7��Ssc��fRV�=�ɣ��!�9� ���9�&�H�<e@?�L�o:e������H��µ���� w��g&L}�.��ф-"c8O��;�z,���h��sB�"�:�(1f�`1e�f��Ä[sR��V !Q6�9v�Sa�sN��P����=�r�F�۸360"f��'�`:��J���� �=K��$������4�:":;4�y�?�9�[ fV����/�^��%�sP��nX�	���+��,�˗��;f���@��Hխ�b�zB��2���˩��#�]�����Ĥ�}l�tܚ�G���{��}s��f���G>�a�B��G�{���|ƕ�׷�I0���$�mry��R�h�	x�J��lE�~Vλ 1@ο"�?�&��n��N����bug=r��X[��i�*]☞�Y1���G��L��ڴ�����O>�������=��7��b��������)?^-YA�1^^2XP�����Q�ÀN��W�1L��s��/��4�\�ݻA=�*��퇗`J[��(p�\Om66M��o,���&Y�� !�J��z��`D�$�!�2�C^����.�X����)�9���_��UO��ya� ��;��^v�S C-� @�!@�����F[ �@��	T�TT�����DG��3U -�a#�r�ɲ���� T��-�U9zB��1�b� ��w �����e7
cD?��r]-X�H*�:�_Z��ႁ^p�jk���伄�ʘ�=hH��ف�� ��9�)�׮8�(J+A�����
v����+�������zFet8*�WfmWh�  D�*��E�� �)��U��#�{D(2��
�{ڗ����uyk0b�Y�䅋C��G;�1Ր��k� ��<�Y/�$�!�7��Wj�RK�|������Wf��]�ʢ�p/�V�x�`�`���5�HVI?��D*��j��!��z1�R�!��}	ۅp F4}����   IDAT��ȵ�fdTc�ry��^�Fw75��;�^|��fLp]Პ���؈�pw	�;j�6=[`3@��*��ȥuwII0{�x� �������oܚ�����C�neEV�!s2Q�R��{��r�uוg��3�G�9c]���[F�}���z��o�V�'��6�<��1�	�A_f c��g���z�-��OQ��Xtm*�ڶL�H��jF�R��n��!�<5*���1a���i�Etx#�U��^��=T�G]懂 ���R[��yJ������E�l��ܦj�]~�wV�)���#6�n-ڰB M)9�0�x*fԙ��EӋ��<��lU4ǔ.�#�٥Wy7n� � ?���v���Z���(E�C��%,~x3Aj'T>fT�����1�H��X�7���N�|LA�����Ź2C�d� �%͈@�%b���n��ϫ>�4��
X��31��}UgЇ;���9S�l`-�/t1$�P�bIg�Mqo� '/ra��]a\&e�ڕ�������(s�.��.�5��V��)��T���R�R�i4[�5�Co�9nڴ��OZ�� ]�I`ڄqI��1��:��=�r�`g�y7*��W5����$�Б��"q��N@���L����H6��*�M�V���H<����R�c�oW�����3��W��6e"C� �k 3�U~��7��|j��<Q(4�5;v&x��^��C&f�I\p��H�5�H�hw����(N+�c ٤��+M���:�MJ��1��pa�6�9?�q����%֣9��(5��`���q� (�sb�`�j�i�	��}=����c�z%�~X�� t@-�l��w��]J�U�n��W�������t��+N@�7�c0��'c\����>mtT�L�$���TG��A����kS�T=�btG���J�g����e��yj�Ij���OM,���j-bɵ�xY�
�K��E�*@��,�;w3���šY�F�A�;QS��y~AeaܿOy~n+�u�(�E��P�w�X�(P�!dmv��2;�V�,U�V���O>E.�=1E���hTK
Cc�g �A���Ls�?�7���QUH!$!�Љs��
c���*C�>��]O(|��a� ��!w��\*A��E�AuX��̈́l+���#�#��� h��4t&n[�l/ ��$zYl�(t<�Fz������b��B�;�\�Ղ�̑7	%V����>�63ЙUԞ .
>�0��;-s�p-'�������꓈`���j�"��7s�[�#�����p��]�� 5��	7i?�����\�Quj+F��r�F��5�| /�4��0KT�Q������)�Me0��Y.����l���{����@��!��Z[p;�!#^�e�
j�>cd�Q ��WtM�7�3_�$��"b�dY�|f�L9��g��.�M8�s3�d�Ft� HZG�;ˀ8����O!h��2ĳ��sTm�L]�w��q)~��D��h����?�Dg¨�Zֿ������� �c��.f�6>KNe,Cbg�����Tʊ6��ڷ3j���S�	��d�O!�׵a�xx8��vɅ78>��\*�*h�
$�+^�_�u�-R�6&�Z��:���e\l�"tv������q�����kA��f�\��esa?�74.��vM,SdC��creQ��u�Xt`г���c��8+�* 
�NMg["��O��R�^��[�k�+�߫Eh���Ұ��=h�u�9稀��f�>��ăJ�ȇ��A~�[:'׶�cgk�1-h�0��@�C$D\��B�6j]�����6���X ���@]�C@�I�&��aq��Q�X8�}b����:�� ���rn��	�<�\) *
�E�)�^�kdHh;fG���j�7Y��?�`?3�*�dd��R`P7b ��\]]h��>��U�dUG�2uR<��G�*v�$���4�e `#��耘r�2�H�QD�ъ�Bn>�3�A�̆���`4��0�#� ����s�|_�W @����>G5�97z1oH�0����{�KLFS-����V&��x�f�)���B�X��G�D<�9�ZN�5���=��,�|F�6�XW,ܶw������y�{N��?�Y�{P��������w ��abn;5�cF�����dA�J��/D��f���{����u�y��p]���B�+��&r��e��AT�;����R��]�g�7�j�w:ˠt�����:�+q���zmJ_"
�+w�A�?T����D�Vvw�9�GA�)#���K����+�vPE�>|%gT��4qm��p�)��@��Y���1���>��䨀��T!¬a�5�t��C�էr����&�Ώ�Ո>��\�~����%�5��X��֯3� �T��������o{AA����'ѲY9Q���^(fT�͊�K%]eր�c�*�B��pW~1�e����W
���CJDYͫ�r,�a�c���M�UBs#���Y��f��h	��]Vƙ"�0S,�Q:� ��6�8\�"�òTwE�؏�&7�Nh 2���F��;�9��DD�XlЂ5�}(�/�~`b��Uf��>c��3|u��ZO,�5���n��*��
`��]:O�Y�	��F�[&C�.2��0H����E5��w�h"b'Jm��2iWe� ��qz9��3ˊ��cB�	��,�;�GbS׃�Ǻ�`�t~�R0K�S��߰-�:�T�h���b^h� ��Ɣ�w����s�έ��;�,Y�����TjT��L��k�z1@����{�,�k��u�P���4T�/A�YT���Wd��te?�3yz�h9j�6� F�8���|�M��S��A �% �ov��� I��c����Iͅ~�����0��d�&!��ilzڴ9SZU�P��߿ҥY~��^~�!g�~����ʐ���t������3XfO<�w�QX XZ+'�p�O�jo&ꆫ]s�����<�S%�n-��8P�$����UR�A�16V^+�v�6�U$E-Tg�⯟�Xd�k��(�4�^D2�p����#ռ&�����s����RP9�p��h2�щlB����p��Y��Q�'D����17& �b�M����hvh��ѰvSc��Y��.����0#����d��n�ܒÆ���;�&+D�c�Xܜ,��A�~���H_�F��04�F��"�J���X��ŁB4	�#r	��H!]�*@Ӏ>B��Z7��ɴXڸUMNFq��#D@�T�
#�9Bۓ!��Vm�����̔tOji mD�0�� Ȇڠ��6�\+�0����`E¥6_c*��0q��<��"�3�^1��O�������Tc0�G��864-�� �/ے�@#�A�����s��xL9�3����>�le�~Fy�C����U?i������T̃|��$t?��C���@�ܟ�j�`��B�7 �v��X���>��H�s��{v� ��EϺc����-:3��x�8�ɂ�
��8s-���v�����Z� �lW^��R���&fs�Ϗ�Ž��e�ÏY<~��&�<�w��9�!�ϱ������:�(��1��h��hk���+�?#GV@�k�G�o"��3?�ĉk��g��qY'�ED�w�����Qf�E����ٷ�������;���u�l��)�o�6_o|���:q���8yS��tp�6 ��LoZ�|�e�����L�a��x=�aXb������8w~���Q�>3���nl�1%�z>�By0��ڧ���V%�ӂG">rgP_jRB�Equi7�����o��"0�]��(�� Ǯ�X6(�F�v\�Z�o��z�v{gժ����B��?FA�\_�x+��	�ɢ�D͠q��i��+� �=.*�S�W�V��G"�(��ϵ1 DFQ*��M�@;<B��u>tA��tYv�Zxq1�y?.���ʈ�CV[:I #J�ȱ����R�&������ �Q��������Y���dd�]�lPB|�g�Sʝ_ù)�}3�>�������B�թ���i�7Qpɮ.�M0.�����W��>�AAה��]�����zֳ~����,b\��w��u���!ȍ��z��8��O��&��n�lG��1C7S7<��TG��P`w�\qI�-0I��}�߸�E8`ڭӍ�g����� �pfu.�gw\F<��������آ�0���>������3�{0u@�����y���n��'� �����%��Ч�b�f����V�*.aAz94��/��Y�k��~�Ck�9�O�������2�3W����H-3_�a�Q�eY���UB�%��-�il��6��P��1m@
֗���kZ��r��c{H!m�Q��� s[�lw�@g�"�(����\�a�"Y�@�M;��9]D�G���6"5FԮc�0W��4��^b���|���{`��k`Nq����@���b�F(F.�C_���[s�t��V"�&_�Bx�|�$��M��ain��cnZ��2	͠ȅ�G���ŤO��֞�t�r�vlDfj��L���)�� �����=u�[P�t�M.�� �*��;��f�%��,S�� 
��_��`���C��CaF-zYu>Y��1��`\P�D��ygN�&Ј����Ε���{\gXf�}14�:�$?���'hS�IjuyY3#k��P-R�a>�)�A�[<Z��v*�Q�� �\��ţ��0�f}%&�ς��"�P���ݔx��i#��(n�d�<O�6܀�­���|r�Ufʺ��J�=/>�9��tuw���v)�����#�OI1o���S`d�4B{��ا�s�
��
Q
�΃ԃ
�-yoЏ1ga��p.ړ�&YϜ����VkV���=�7P{0R2�
6�l���n* �Ne!87mc|<_*���������]&���\6 0}�{0Fzܰ�A�����}Ŀ*�K�i������K<O�����[���Rq����sM�z~��YtA�o4a�Hh��F�繃:G�;< �ni�@�P$U�zFѤ������y�7��DGح�oʬ0����QE�H�P��ܪ5���*��D�_�jj"�Q��ŵVe5V(G���Q��K\>*P�u�H:ʆ�/��/����7�+[��i��%߽����o�{Ri֯�:�M�XO��i��W�C����*�a�ܤ�aQ}v�����1- A�e�� -��� �v~7��hr�]j��3z�[Z���%!����Eƿ�#L2)� �uƴS�P��
hav��ܖk1�x�á��	�C+��P�
�w�$�h+��VX�a+X�X �QHS��I��|x�f �Sp D�2�J�n ���)��^�2�.����<�!F��;zYӣv��.ڋ� ��v�2�b}l�|�X��F�9ޠe�����6���S���8C��vH/T�C�R���'��5�@�u2:!���]dc�v��v#�R����W��V@�q�0�w=2�����K�M5p�u,�Uw	}�c<N:�de�]Qv��D����]|��v?Ў�ڑu�	�� c0y�P3�O�bi�Z����4� ��(���/�G��e��p�Et!�������-���i�) �{>T&	pD3}ܾvӆ��� ���{jk��h,�1�m�S���(8�+��s��]������'�#}���XF�`P�%�\�VnB�c\��0��i��&ɜ���(L�$S(�n����9ah}F)�C9�K�tTnz��s�A\�����q�K���,]��c��1\��F�"��S��q�>p����׿Z�UY��N;�l���T��%�sܹ���i��^�U���O���L�a�q�5��� E9��ٛr�vd��§�"3k,����-������x7It�Q*�w��%&C;+�o&�9a0��D5ô`Hud��9�X�z%T�i/w���we��~ة�q����)@C��Ek�Q�0 �s$���8"Q5��Е�!A!��@N��j�$����ذ�"^�%�r�Ο���~5�DSm�"���5��zA��1pVae�G'��)�$?�#�H��@*�^�:� ���Hq��pof�zlӳ�Ny�r�]��iGc���d�0Zb�� ��
�ŘQ��A�<'l�j�=���l�LP9'����f9S��	��5D�q"b�\;M�י�f����nL�<"�&�t�:A���fX�2�Y�9�h�6B�q�!$W��.H���V�l�����0ٖԝ��rm.�O�ie��N@)Z�Y�ҍ�&���!A��鈢�3�A�L-�j�+H�K ��� s�9�9�kOc��G��(?�ju'1ޞ�l"
�MTٚ�g��-D��Cn
��� �|��7� ��,��q����.���l^���*�F��1�ٲl�
�A�td���SD��t0��g�Dmt�I��XJ1�&���k#�W�r�맽m�#M��`&���k��}��R^��=_p�M�h}p��&r�0�~���%�������YH��]�J����ig�����+����v�ª�h^ZK��pZ�V�H���a؊ů���E&�0�F��)[f�O�燩i�y�#�8~��3��E�B-����4�;X��y�aт]�8Y��!�E�L�^%�;���S�-��z=y����%�G�U%|J(�(�)e�V��q��9-�,�$-���c�,7�~��ګ쪚�a��Mq���ʡ3*�t��˪�8����C����ۨ[c�����;..m�\���~�G$� ��(2@��( j`��(į�J�\2M�H�@6�ӂG��nh4?`Q��2��ԧt #�UvY�!M�DٷG�?���M(d<ht��"�,�unZ蝹�z�wg�� �@�v�wы �e7�O���@?�B;y�t�l�1�'��L�5\�������%�:ҏQ�+`-�#�*s�DԺ�i�S�ש����<4c���n[�'��v�C6t��k\3�i�	�+D��oGQ�ڙ�M=*�:)f���9�+�U� cءy1�Q�n��Ʋ�e�-�b]��"�0���,�Mt8bdGj&��Y��"�
(Q���p�.�9���'�v
�G���sűT6Oc�k ��ѩ�J[�9�v��<L@�����^�Q���%U*kn)��`��fʣ*Κ��'z�ρ3��(g���]?N����O���eY�̺����$e|u�V��c���p2ʇ�Ϙ���B�iPX��SJUt)��ʜ�ɉ,%$G�?���hS[ft!^̥p�(#���J��C��5Qɞ�1�?�3{����h���m�:u`�6�"����J��m��l��2��5��'@:�cg4���!��Y [[7ͭ����|�\u�b�����_�6cZ;�` (km��_��Y����"tCV��E@���?�U0UmKLK��;6N��#_�C�r�U?P�5���~�g	mfW�,�+���G�0���"����
p�����Z '�e�t��n�#�Ԃr��7�uJ*�y�rb˦ҹTQC��3��j���阘����K:X��]��!ؙ��c
�5Ô���Z$���J���~"�0Y�#�lZ����!J�~��+�r���iX߹��ۜ�xRmb�O
5�+���:"a0�>oU��
��a�yj-MK/��|���$Qi�y8F��mD-���o��5�G4�!�˱*.�<�.�ta��m"W���2ڴ���:�0����M��sN"�y�R��GT�D��n���@�N���� V`킄�r�^���p�`�Cfw������b`���΃��o��C��}2�d�$ÈA�~����w�v���2�����$%�c�G:_��sϹA �	p�n�f樒.��� 0Y\���e����؍�)"qxչf�,�� T��b
R��V��0����"�>�aD]�T��}f� �75�-܄o������=�F`z(ܘ��� 70��bԩs�c��)� E����1"!b���#�$��fb�?'��6�a�**l�u~�tJ�]֯f�Y�X�)G�+�B��Y	��~��)(�"�̳�<��q����5�;�s�u�63\K��`�d��%�p�;E�zLl�n@{�Y?�_��j^Sό�%A��V#p`�D��s&n͉�Q����R?K�D����W6)O�*�ؤ��ގ �M��B�wsm���(h~%���c�	:�1�3#;y����W��`��Q�O���7z�ͺ ��]
A%[-�r���~�������}2R}�\Љs�9����ZDHH�S��]8:%Hm/va��٨v�-Zغ�1jo��Of'�5���c�pQ�R��	W
����h6�� �R!D4$�cwR��ZA��'�oF}
r]2��q�m�U�Ͳ蜔1��i�\d�-΄u��w�[��1�\����PV�n�͆���2l�!���C��mAj��e���F�s��`��ϺG�H�?`� u^q5���9��K�>Ǖ�¡�J̙�Kb��7��Z^vu9^Cc�t
_��YֿRI�-~��r���hǽB�O1FU�ù87�����Uv#���Q�*���^���hG�D�	�F����ŋc�$���7�ol��/�����4�8'ғq�ֲ�o��׫,�$�L�0hjeUw>�oS��: ��L�yO�$Μ?���炙+��6��q��w�¬ߕ�t�'��o��a���8�tK�� Y���f�D�	�����2�ų�3�s1�VZ�铑�9��r��Mб�]����7��-�ɑ�~�j����y�`N@��qk	lV��2�Z7XwAX��[��U�ݴ��a%�lW(�D�P�sb���P�VT�'��7a�gt�ܖ���ƤGnᙩQ�h�V��Ea�K?I�/2A�9��_����B{����c4�@?\��b�w��6��8��&����v�h2��[�c0<c#���|����q�������.D�*1�*��ev(�<�m2�=�ϙ*kǏDQ����NeO��!�Ɯ� ��ؑ�1�Ckbwn��(�Y:���	$�c�ć��!��.��n)D�S���`���Ϙ�b���kW{!&Q����H���е �Z�b`�I����ar���6�3vd��+i��7̂� $�7bC���V���^h�Bf#�P�0İY�*�>���@PlND�D��S<�� �=Mh������P�fڕ ���Q?��q=-�3FCͱ�/m4�P8� 6�2�YS��ͰX�O|�S2t�˙g��q�`]�F�Nن>���_���__��A�KD^��y�J`\���Y$.`ˏ50���lT�K�1O(����)F�c�`~������ �1�.�u�p�dɌ��m�=�����`3�#�ŋc�K	x������fD���/!��l�*��|��
�׮B=���	�b�G!Z�3�!��������f���g��V��
��=d~,�h�c��	�0����M�RIV�ڼY�;����;����kw,2'{%wW;ωj}�/W��и���ݽ{�ֺA1A�c	 զhQ���>fX���k��}7��Gsp\�3&'��5�m�f(`�����LA*!_��fz���ô�?N__A�1Zf��Ө��;��!��Y����.���d���`E0������� ||
q/>{��T�&tW �?�y��=Щ�1�z�c��\+K���zbRt��9LRE!����{q�`gE$E
���aXj9f^K%�D�aw@	V�
NG��&��Ν;j�
n�������85�k\<�d��AY*&��0`���P\���4BZ�%6(�@�f��U��f����axj���z�[�b\޳b�M�{�mF���B�@�����d����f�N��$YG8�C2���O�+������t.�U�Q���w7m:� j����O��Qd�>��m��r�^hI���Hc���b@с�������v�3��_?��5;ˉ'��H��va�����_P.���EJ��d�0� (���(ے��1��6�$�\x(sܦf`����F0����� ~�H���W���g]��B>�f;��2��(E�W�l�D�)�yN6���^�J���Pdr���X��8�0���SG��:^v[R)����xڗ��X��AU|��x��x���/�LF0�d��O�!^v���s3��֘O5����� ��iLp�nX��������v߶us$U���L�p�w�֛#�?AA�r�o���mykY&`�k�N�X>;wl0"g�)�	F����C!�Z/n���#�;�t��*�PE���M�UǬך��K;��ZF�g�^Z�ha�-����� �0F��@̻��U���pe��ra�nd�~D�LQ��ع�aU8�w�,��4f%6���tT�a��$N9�$�49d�����1-ڰA��Ds�o(�t�	acH�?�4�-�u�^M�E���������H{���E��5F7��Q���lD*����k���(^ ����Ȫ���8��r�"=n���؝�;�fi��C�Kc �DY�m:`W�V�?��0$�hX�A|�E`���l�F1� X�FM��-��LP����3:#��t�ѩn��=�
���a�aÅ[�蜚Lcc������ ��A�v$� ���[т�v����c���0IR��40�N���H;}w�2�M �����@����2 @s�1G� ���6�%������ng� �x�%�:�&��Am�~1������S�=.�v�İ�蚍N�h��g(�*�G�j��6�5����'��s5A(׶��n�p�;����`'��c��t���PS���<uT�"�)�Xe�d���A��s�l��Ǽ�儕�5�8��)� *���R�d��zew�څ�'A9}i$���c'X{�C�ļa$r^�Z�������T�cWy�~�ERٶL�5B�Ӷ��,��~q��ݿ�ŠI2J1f�W딈� ڷ�?����b��G�ZE1�Kz`\;˩*�A$�)�?�P�m��i��P�}p/Y#���5�G.i-Ǯ��9�w��������1�R2Z�p�I-��2�����I��6v��H�\�x�d����3���f�hڑ:�X˔4+��yZk=h���mo�)�16�JTeG�-�Z|=�XA���=1*]����c�z/��K�g irw�;��|jw;�C��T��z$VHB(��+�biƴ�_����vl���A��أůM�m]F�A�G���"�:�g��:�����xr�6(X�K
v��� *��`!"�pDu��TE�1^,���p��0�G�t-\$��A���f��CFXt���p������]e��E6��G�#����/Ԧ"��s�P�^�:$'~� ���b`�:)��7	���"�j"�`b)��u�L��1�zd�%��#<�e#Su?K����n0|��.�6}�����~w�fԚ�k$�^m��F&�>1��lOʴ��O����=.�V��ރU=�#�M��NY�!�0"��D�B��;!󸬔jA�s���P;T+����|���g?cƈ]��@nT�(���f��<��d����H��A��F�FȆ��S�Ǧc�4ޅ���'�H���0�0S0-��z�=����?�S��_��Ѱ]Q��=���>�	>b�N��%v�Sj���\2/`�h��`#�F��Zs��0w]?�nu��V�9�?��V�<Rޘ��lD"�/N�~$� �2����j���J�ϊ�JPB��W}v��7x.;i�j�Q��<@S���scT�a�'�Q{f��8֪	=�۴6�yםe�j">���]�Їx�B�i��ε���厛n�i�\\Z.W���e1���%�	�����*�k>v����t��������w������+���O6�v�i�seF�	���l�(�/�mr�wv�	,�"�mY�'T�ar��XAr���4>��&̓f~���Y>���Gσ�x�]c�c�g���{��}��o�����֭�d^����� �~u��Ul?	����#b�Ch}Z�%�����
��)�a���������
W/ǠePv�Q�c��=ZHY��g�zQT�o���`��!!�a�٘�*\S�pSC��#ZN�-��i�/f@~y"� V�(Wr3Sn�sk�Ff���~��s�30 ���9կ[��«bf2��{�1�1!�U��Y�M��m��b���A[%��~�p�e�9�pBٲ9�P��!D�AQe�]��KE�R8?��2��"3!p3.� �B�Y�S�M���4Q�ÌX�1 aͬ��B����r!V]?��Q��R��z�Ȯ�B��Ex����,.y�ZPyU���]96�D��0$��o� `�r�`��A#����NY�% ���� ���q��N���`�y�8 5]3~����`e!�yIC���V�]��KU����>Q޲Q$�E�����E��C�Ir��W�Y�]M sZڝe8\�������k��I-�󽸿��u�M��Zus�A�6Kj�(Λz�dar�Hp���\K���������;�eo�<j~iMp��3��6����q�Yֹ������i��u��Rx�`a�5��gրSN9�<��/�w��U\�c=��m[��%dr�W?j��������v�˹��;�,�.mH!��zV>RRPv���=�ts9r��r��e׶���պ{�{�FĊ��,K�Ԭ���=hfp����c�h����ޣ'��7�L�U��Y=�3��Csʍ�����*Ay3�Lx���G�,D�KӐ{5�cѤy֤1֣��$���ޜ����={����Ϫ_��w )~�f�,I�65~��'m�z>�l�_8��f&����>��"��]u��\/z�S,�7ҷߎ�	��B�O#͟W�$o�z���C�ª�	B93�;�,%�Wj+%ج��>�� ��-��"*p�,�"3SA����uN�6Rj{*+�ع��_�����2���Xpt�R-�i���f��1��f�,��z�����[,�D�X�����YaW��1I���Bx����$��}��� �FQ�@�o�����^�牭@ŉu����|�
�=����BM�v��lw�r!�}��P�`" ��11�6�Du�1BN��� T����'�e��$�~YЭ��^s�ϕ�GqU��2�`!Gƿ�E�P��M���.�9�׀ň���;Ŀّ�&'�����R�D���ۣb�0�g���/���̂�-R$��c��]��H1q>\;ˢ����e?A	2+�r������FC (uX�^����0@�1���C���&56��ʟD���\k�v�k�7B1�	�l����&�~��Sl�\�lB�>}�k�Pju!�Ʃ����P����5`�{���}�K�Sܢl|�'�և$������։�p�`���7�0�r��R��ti�_��ؠy���� j����G�
0��}���O)+=v@i��ե���NI����σ "���=��rm*_�2cM_H��d����K�W���Q�|����="�}w�"#�X`����y�⒋ڛ�g&2�r��֞��&1�M]��M�+�^��ѓ�4{��=8�wL ͏3��pe�9��p�)������G�L��#[��FS5��_/�����f桞�qM�s���J����qۭ�/���(���g��u�f���/����a��/�C��t3���|�&��\��F��ޚc���F��{�`�Y�u�A�6еt�YQ�����:�墎@TWg!.\52f$�`���.}����(a��u�)\��+n\/,�s�Y	�'��s*H#) P���.��[jw0���B?אav�XO��'g�K�8��4B/���}�'���X`�ѽ �F�3�E�.�<D�D�9�cT�m�FF��-bp!C�^(\�c�Y?��Tʂ�:.h�n֒�~�J=����J
��!�r����.���X3WN��3��1�;�bX1Xb��Y6�G��5����D�״��%1n* n.j�9�Jk���LW5��/��a|q��( Ee}��c�x�`7"�Hԧ��*��ME����p���ۈ�ͱC7������y�Դ�{��(ߒ�X5�O�p#s�n�6y��K�K�r�{�m�λȜ5����j;��b��n#���4�bt�����I-Tc!�!';�s�g�kTc�yl����U�]�I������ Hce��ƀ��������r��m�hǈX��{:'�"Ƙ��X#��n $�6z�	��� ���?��'	�<�"v�g��-w�&��z
��C[����+&Y� ֨\����9�bgר�R�!ˀ�9��(�P�d�t�4u�@U���_�H���%�*��'��Si���9�3���:��έ���ۮ�٥�V�k��Sv�I���MN���ܵ�u��AaE]��)L� ���.lV}������B����:�c:^�j����푘�q=�Sz�E�D^�0�@�yi���;F����~}w1��=-�|g��.�o� �maG�'=}d��}�5�Q���6�7��ޮ�e6���L��
U�d��UB�̭Z�z��wꁇ�=��	n1�Z��5Ǳ�ڙ�j1bW�}Xa���԰U��={mb��r�E~xv���홁"���퓗�<gb72���� ��z*���"�3N\';�q�lk9�\1��`��$������N>k+�ǎH��������a�N�a'�Ӡe��Ha4���o�v�<��Q�� q�
����oټ��`B�/.���93\O�E�#���)�5�S��`��C�		L���i��2X܇� i	*���Ǚ�TB����@;>cl�MCBԣh�+C�D~�Pr�(�6�1!��=C�����K�6��+C�>8�5�T��f3� ��lP���lq4nf����_�T���p�nC��
���6�Oj��d�0ܩ�q��\�w��$��ݩ��ڎ����01 ��`�]�{x.�������nV�}Οs#�,E�K� �1�q�<E0�� 7�	2��W/����-2�G���B�|_��7'j/�6H�� ��{N�����au3 H����sJ�Jn(x� H����n\w�u�r9N5�X3wn��4}(�n���\)�Ї��J�z����2>]e�r�9�h�z�X-���;��N�/����v�TT\�+�������=�����ԧ����
�Ö���3E����+����7I�<973���;��ؽkjnJ��-sJ͡�unJ����a\hf���gi���&����I����Lͨ/g J9_�r�j����������֏�j�����o�����9a�ZE�k�$�W���6���X|ݯXA����~06[p>�L/$$C�������].@(��=�P�} y@��s�ߴ3�eJ-��ј@�`"@!��,�$�Nh�&wZ���+�ɕ�_c����q��[sd٥R#2J���r��
dAC{���l烵Ц�2���0�m�ŝ]L�o6Վ�F>B����#�}�_�����dOfv�9%E�А
�R40�	Q~ ؎�Y	��b������ט�H9�Ō�W��Ϊ�W�-P�����-��e�M�?I�a� ��0Ҥ�m���x��٭51"Q6%
Fm�ۅ{1��Q�o�k�K_S�=��,��� I�/,�+�{�[_�83'�YƽKF��3�x���#r�!�U�^�~��JȺݮ�*�~�x�T���D���1�0��)!:�������Y@�P��p#��9�Lח�ߐ�j�H��Y����g�* ����w�սH f\��_�9�>s�~E�߭�c%v��;D��{�Q�CT�^������ʫ��G� �'�`���� ���d���@HX���7솎c~����T`�L4��cC����1��殻'�c�����q���zp��6か
�>����q�2��]��M��ǅ���.Q%�J�m
9g�F�C���w�Q��r��ǔ����9��E����g�"
/����ȇ?̌���|���\����5�����u޲m�J���1�u�Mײ���s��A�o�jW\7Qg}+�	ýLAc�U��nrwu�M<἟Y��'������,<4��$��":��S>����fB1:а9� �)�
4��Ր���~Q]]#���q�b�a�Ij����:�~,H����
�1� ���u1��B�;jn}L��2-�r�Ѧ&��E��vO_iV��Z�Ě��TVˈ�|�lA��sfL_Yx]hSL��3�mj�A��Ȁ�9�+�	�O�vU����u���I-XD�E]'j*!vh��D]+��V�}ø�q���(�5,����]�!#�Ga�,�d�&�G�#A���V������t�,��RV�l������ʡ�Ӹ�^ppզz��p[-ފ�!���&Ѓ�i��A-��qR�^�@LYgF��`ȴ�ӏ\5���|� *��%6Z�kN�^�H�[Q��lR��4�}��ic��(T�%*QQN��Ui�=�ZT\��0�  �*���;lZ8�I��
t8t(�]�� �»���C�NX׬Y��
�Rd$%DՏ@�����A�&�W�~&f�E-�UUH�&%����xRbě��41�S$z��ʳ1*���KpB��!'�=�n�~|��������Ăp�ԝ�I)`�S���6�H��:a�HE�KʸØ)���A��u݇Kd�H�; p�x�Rp���\�t\�,���g�t-�U�m��~��z���l�K�賌R$�r��o�И!�Í�����E�1m::�ĭ�`C=;�	�]�vX)7��ğu���+�+�W~��5ɥ@5�t�i�]�$���zr�S��q����&���oH��Q�Q�'�Y+0:��6���|Q��6+}��q�'��=JܸO)%��?�׊��|߫2+������Xq����>sfa�?f=��c�`�����0vQ怄�5ח_w�D"�Ljb�������kMGDJ�Gi�)����M\�n�a�N��:�DD��'�/v�Ӕ�Htu�_���9�\0EW,��n�^�@����Yg��Zv�~k^B���O9�!�VL	�����������3,�2 z��MU�.1�� `<�����ȒL��
�߸�|@�̌��9�c ���E8j������]�ڟ��G>�����C�=h?F��	�� 1_V��>�Q�Z�ЖK{aם�qGya����Z��@�{H����t�߰CZ��2�P�#���Wax��& �5A$�Xq�Ї��1"�����g4Rf���
E�	Ɩݻ�zڭY�GQ(Ww�"���N�dR�#3sɂE(��EF4�I|02�P_����_]`��o�Y��RG8�b���`��U_9c��F�!�$���EuUq���{��%���E��WIW?X�ԉٍˆ�^;�,��byX�5��(:*�7�6D'���(��� �\�Mmh�6q���l\[|ϕ\p��&
���7�G�/���2�\��]��s���I�s��y��#�<�d��*��sr̅��۔;�_�zy�c'O]2%�F	���=��~M9Qn3���A�(��:\����l��������ԍs���wͳ^�Kl�Z׺tyYջ��a]����~�Fk��Vj�[������ڴ�(�G؝���A�a��>o.������:_��`-���O���K�Ԩݸ����{6�6(bL�v(�ho�arp� �D״Kǔ_�{��`d+F��/F%� ��xY �s`$Fw�28:b�F�\2�-b�L���.WH*�3��	�ЧqC�Q82�W�E��^~|'��oY���� �ES��i���}A�햱�z�V*�M��.-�,��p
�-[��]L��1��R���H`��؀\��j�wؘ %��������~ZY�Vn �-b��  /e��D��ukו�����F��U
9'pH��h�uN��܊�:���Y�	�	�3��X�aX�$A�C�RM�5�W+��6��$EH�q�ܮ����'@^�fK���lW�p���� v�G����-P�AtD�\���t	q�4M�lٲ�Y�!��=Dy�`�l�a��7fNqU����(�q��,��������"�4 $bޜ�hY�)�1	�8��B�s��:i���2z>ȭcM.��}�縌��hb���G)�|�]�'�t�57��O����7�G{�8W�����z)VOV�k��Eغu@zq�s�y�Hj^g�!�v�]E���'=ɹ�`u�%�&�'?����}�s3B�^��NP�O#��vn�J�0��y�c�Z��CNi���	�X�Ʋ\�7�>�hi�FU��*/�p����5��s�v�_��aΝ�Z�@th��>�&6isb�F�r6��CG�蔫�˕(�p����C{*�Y������������":���0��� �&�ҹC�Q�0a4�`�{a��`PhVh$���h���g#;������jË� ����b�NI�(�H�^,"Z�v���z��N9�e(�,�L
,��+{��R�
_��\��ػgo���z��"���oVE��N���)2;���4v���i�^�pQ]�u̴��v%��8l	��Z��KeX�1N�j߰n�����fu����`Y��;`����wA땺�F��]:G�y@L�.19�(Wʄ���=���˥�^"�q�r�l��a���%C�>%��6k/8 n����]��'�- 7�d�#�7eIb�)� |���"@��"^E�Q��?�A���?g]F���^1Ǔ}��T��cN�D��<ĺv[yΔ�n��|�_,����A�~�ܮ�����+��a������fƷ�A���̂�+�3^�:EZ \Dοd�� Ap�@��O|�Jhy����^6K���c��?��r��T��ps3��ݬ8�[�·���ߩuJ��<�/�^F�e�E�
ox����k�i����v��/��G�N�� I&��s&�I�'�w�K���s��O��f�*�F;H~�3˜��۽|��_��_����s~ٺm����g�ē�v�aa�z��`� (h�8n��-c�$�6�.�d��{+Uje�uڨ(7�zs٣5g��b,��y-�94�[�}�=I�Dz�a) OWeOO�<H�����vP+n;�oFa�d\_�D	�3�6���G��Y����=����M%�I!,��tdT��C���x%�t(����cTS�T�ֺ�蛵p�x� B�(M~xP����~Ƞ
���W�\CcZ�����@a D%r�m!+@P�&�KK�dN�׾����x��y��>�h�O~��(�'pСE�Ą�s\��;W��6�$�]Q\F�@���>�	��E?�x�"�F�W@�ý�����]P6m�Tr�C�7ܨv�6��я~�|�ӟu���64(�@��e�=���Q0SQ#A�B�x&��q%��J��+����YgA�$���הo�;����.�[�6+Ae��D��Bb�l,��a�vb�I�X��:ܰ�Ox�C�p���y��(/��x�.pّ����q��j��s��\y�{�+Q�v�t�%��\(cya�+jӹ"��K��(��Yើb.� q>�э���i��_��r�"������|�;˷��-�܇�)ǞR�:묪�R&��t!��Q��p�|��B=1sF�N�ӣ�>��$#�n���}��o�+����=���ɟ�s�{t��W�^>��U���o��\n��k��`^Υ�a>�� �d�8ֆ��¨�������o*�{��̚|�0� ��Y�����5O���@��	�
�D�_\Չ��P�y��׈�c��|�����|��Y.���b}>�����_(^|I�� !�s�4>�@�mĦDz)�>K5��EF�P����ފħk��c��i�ֺp��7I4���Yܵ���E	��*�=�vz>�~F�'�>�OaZ#�W�A)�G ����r=��dL������&�{��w}rC��̪/�ǡ�~�z���OF,���G-d�dy�YXT�25��(�A������Ac?�Y�0��z`��<W��֪��L� ���x�a��%cW��(����;��ۋ��c��M��}�-�Eь��f����ɚf�3�(\ﱳ���>�Ϟ�+�RViW7������{G�¬�N�?t3vi�v��L��Mh��*���q�л`lm���Q��;E��� ���/��\tمe�c�O�'=�g�㽫����)�������J"<9Jg�� h��s���>����?�:�s���} ���W�,檩���b����~����o.��r�2�����>�<�ϔ� �����W�0�E��Sb�N���8�7�Xd�V���y��p�J�N$�E]T���>*���c��6������� P����>��t�D��p�Ŝ
=�ua�IP���h`�4�� N�[�9��L����*���»��.�3�:���MZ.���2:3R��x�����=��h&�mDv!��#`�yp�3�׬��_���9R�q3Sl�c���-oy�ٯo����o,�|�9���//_��r±�;�h�X
'� �]�Y��dGV�ŸD2�2_`��|>V�X�/���z	�/��²{��r�
�����q��%%�
�;�|���%��N�Y���$"8+@��H�2�M�ܴ=���sIʉ�E������|�_q:4i�T��y��}��5��	6#]����o`����:n��W�Ĉ���S�y��̒��:a�fs�D�%~�siwf�(��2��U�N8�2�,�o�Ԧ�U� ��@�d1���Zs�Y�>ǂ���)�Et��E}F���S\.D+�?-���$�3X2���Wh)j��y��|��j`4'Iag���G$Z_)��|�B�ךw��|�h�FW�ő:�^ #�� 0�����X���v!�۵��%$=u>��0Z�����1T�޶m�w��׭+�>�Q��o}���W#ˮ�Ӟ���{/�]-����P�~ja������5Qf����sF-jb!��q챻5���\�4��З���r嵗����m�*�-�)$�?�6�+V��� �4Bڳ�C�V#�n�
T�'��t��>��{��q��»\yQ���/;���3�(_��ʍ��X��������/��8U���W*��܏����-Q�Q��@�evC?�n�4������������Շ���T��'>�	�ÊR�lذa^��C�n���`���p��7ㅻmF9��ah~��'�\F�b�)�p��������90t�Vm*/|������Z�K*��� �3�����A��5L�X�t�)¨2�¯v���tDy�K^b��[�EW|�lZst������聲G./X=
�f�-Ν0�"�_ͣ�  ���o�Cߥ��.�Z��t��@�s��g�ּ9�s������%D����p�&�.GRD��s �֯��Nm��3���'������ek��#��-�� 
n�g�E��O�W&���t����]2㙿�Lύ�r�1q#�U�h��-��pR��w)�{@c�};���)��<�X�?e=m���|=�w^P���O+���i\�����y�Ѧ)8�[�<=l$t�ZFHr� w��+��?N=��s���(1V�>�y�"2��Bñ ��
���F��7"ن\�,�$���h8j���H4~�0�hm��ūߏ>�L)�\}��XY�fU9�Me�Ļ���j�Y?�0s�=�Q����+_i0�[��L��򗿬<뙿&�i\�k3jwIƛ�<`,-���87�KU�k�:dkn&����ҭ�Q�-n�׾���6�ַ��r�uז��#W���!��{v��zY��%�J���+V�Qw��zP���u�+��h�P�
�K�V��w�m9�r���_*/}�KZ~�U׸H)������@,3̈́0<j�����D�!M`�;}��n���a��o������ovx9���J�.���lF�x$ӕzG	��Ꚑ�(�T��yE���fH�� ��s�u@J�G��g�g��g?�.J)�v�Z�9	q:�=?�*�k��e������a�O��3��m��~���屏;_���o��mxO;����W��\�2���n�A0@�`���"{�y#���?la�Sxm�����YC�t�a����'�׽�u������g YƈW���:Q�=Ϡ#�"��8�"�^��툣�>�y�s�� `���������|�|����&[��N���Qr,����!�223b���*#�m����f�����кW'c���x¬c#}���B��2e�?��1��~��Տ�����-��vq��"��](��FVYm�4S�70B-�h����,S&i6�c1X6.Zx�������XA�7X�0;)M
ތ�v�z@CC�����1�����)wL�4��ra�A���P���C��gA�-`aA�!�<�O���'��c�._����������� �T#ڭ�u��]U���ᢘ��Jų�+�����׾�<�)O)��r�v���EB�5`�ڤ���Vi�F�f�$p�!�J�D������O�)�B�۶�Gi7��?z��Q_}�U���?J;�9plV��i�ltL�L�4���թ���e' 2#��L?�+ƵO;ߓN<Q��A����<�)�U�z�uS��}B{Ө���ŬScU]f��b8�_�=�[�7ƕW����;��y�'&���7�����L���N)�5\�>�e���Q����f���
� �t4#�~㪠>bQ#��`��@�r�<��/O����k��N�㖲jժ`��W��2�!�1��Kw%�]�js��H����I�.F�?�ؾ�i���)�́���e���H����<|�1�k�U��������g��J�� �{�_������8��V���W�O��dܸЮ�$5Kk��_�j�]��F���
Q�\���$mUd܀�9�5֮�E��k��*t<v�Ƌ�y���eG� ���Wq��|�@Q�"�D�j��$�ޠT�5����r�r6FN��} �b-��Ԉk���v���K�{Q٪����m$�Zy�z�t���Kz��c��]�'����j���XA���bLv�ս��,-RH�Z "��������@��?�i7��S�4o�ݔ
0`sXib��ѥEN�,�{�;˙g�!�+�\��;�nw.
�N)�N���FgU��]��c���n�ŋP�G?���m��#�X|qP�#�8�l�r�Ԛ�Hݡ�~"�������
����V��b5%��
N�>L��E�P�nz���v�a��u���E1 �}ܞ��%�a<#<�b�V@Ye��wF��C�uP�����c�H�~�`a=�łq�|-aX�X\cA�i��`�^X�4���䈢���>�*���o|î�
��B�:�0��`gޝꢛ��<4ڜ���� ��U�v��ۑ���`<��J(H߂ȗ~�I�1����ZD�NnT��k�(s3�3�,�w}�P�y��n��R�Esf���	�a>r�5�\:r��r�^f!2lz����|����9*��>+ǜ���߇������8�h�F�q��\�Թ�ݵ��b�����}���Y����D�)W���с���h�����W�!� (j&R�-`j�6�ʚԓ��H?��<�7)��ǟ����6ou�V���+��Y��kV�&�U,�˒�J��{D��{�z��?�.ߓ�Ɍ���08��j? K���� %���N~�Q�]����_���1ю>��ث���k7�#֮.�ܹ����nk�.N�hmU$�zp<Z[D7.��=J^� ��ڔ�+��C�Wc��;����+#�E��s���hG�����������;v��Uu��ԏ�J�to��7�w+�GG9��ːč�e�B�^'�d��9Y�O���sb���[&������8�@p��p�R4h������O�t5mc�Hُu#s2e( .��`�G���\SEZD�#��T훝��yPٽcgy���Q���z'r��&����Z�T\J�p�e���˖�{��	��;��py5�2d2B3��
�t����?B������nAeܽ�?.P��U�7�7�M9��f�ʈՙ�������O�!�/��@`|0�����.-��a����~��}U�!��V�5�& C�SW�n9������#<\��8�0@�>a�M�)�F��0C�b7���b��&a����5T��7��+��m���r�n�D��Y@;�̾�� ��9�����x�)������-�@�|���U>�W����;�<�ɟf��>�r�񱰙�lxl ��s���^��Gc��Lf�IkwԞ=J%���E/�}��� ��HGs��7������Lb���6Z+��D�r>e�p�M��Q	�a]���0�$���d�fܡR-Ѕ~��%n엾���Q�>�����.���g�>lg4@�j!���R"g�ϥ����9X{���r�D�9�\��&@�`��q__�L���R6o�Vz$�n����C��X�^v
��:"ti�W["/$���L�����WJ����7�������τȫ/	 [|���":��FX"��=D�h�70�.�0
���߬v~$�?Oc��c��,���F��<�.�C:{Xv���O+�=�Vt/^����N���q�-�v-�hH��ޮ������qS��KY]��/eFm�Q�UsRHD��7e΀[���*��J�`)ιC��n)�ַ�?��?�����w}@: ���N@��?R�"��DEA��\@L�hY�]��N���������WJ�i��3%L��׾�E�.���f�5Y�^%�C\:�H(J�ȅC����WA�{�\1���
 �O �����ay@��G�������Z.a���o�^���~��ڟ��g���R�����t�2*������
1O`G ���W�A]�DY_�#0�j����|�ϕ݃��	G�P~�E/*��0�[F�+_���P�@����b��`���	E�����NJ�k�r��:@����P�åyC�D�Q��8�fI�������S��d���_�z�K^�1�-��w�y������6l�j�v�b���B�|,A�1.O@9�R��Pz�Y�?�hū���T����|�3�g���7����;nuH�Źz�)�k���'��a�=�@��	 ��`��S��C�����o���t���e/~i�9�������hJ\�_�җ�7�PN�p�F���u�^c��Z!��Ө ~�� Ak7�9�ŝ�Åf��n�Hv�M�^0^��V�C�X�}�k�y�=߮�W����VQʀo�������E?�ݙ���P3�5�������])�s[������������������4S�G�K׈��\��q}�8�7�ֲ�@t�۾��p���ʋW���r�� �6��ԓJ<׳0�*
�s��y�a%����A�a���Gs��)�Pw~<�a�Q�;��7]S��
�x��ӭ�,w���N�:dG� �f�%t�(e�%�=u�x�_��'�jG�����;.��k	���NHfbbT�e�s�q��c6���S�i�>�B���(_a���
��� )UҴ>1@�U�pǎ��L�_�������?Ӯ�k��/UD�[�t�)'�e����˺Z�.�S+�+����r��LJ5�U�b`���Nѡ�h$F���?p�~�#~�C�+^���'<�|Y����u�/w��p��?$*����EB��q��&��RV/�h`�X�c(\`�p� ����ժ�m۹�,ʳ��[��������c ���߉���w����o�v���m�������˺�X����<?��0v1�j�ժ�Q��믻���#�ź��g�f�%E��^�Gv;|�;߱��Z%�2a	���Q|�+��`�\��/ ڬ��ss2�v�B�d �Ec1VKpt�ڧ� D����g���e��!	䟾�O�^\rɥ��\v��N���I�� �� �w R�ƜhBv�/Q.& �7$�������a�TDխ���?�1��/{�4Q�ʕW\��I��?x��������m ֗a�()ӯ�~�-��<rn1vu������jT# 
��l������C�:[����D>��϶�mo{��Z�	�spۭ���֊�"8FS�gk7$�`	��L ��{�3�j[�k��S㣠��0D�����E���V��;R��8��.�`<��qJ�Ԃ�0K��$�&7}r睛='tփ4Ǘ��%���`m984(09��P�s�r�qh�hC�9�rg�ah���Iz�� {�uM j��m�����+��Gʵ��Y2�kc7�����9�&)3�>/���� �0�O_�p�F�����̀
�A�N�{�[�M3��3���f排��ˢ�?�E�[o�N=�+��`, �U�:�zV���as$�X�~eq�$z�ݼ�B�)�`#4W0\vQ�����s�G<��7~�Y�x�p�1��/����o}K��eҥ��3ɦ�s�b8�X��.�;Ys�y�h3�E�$��]G�E��uQ2���4�v"��:�(�-g?��J�xC9��W)r��22�wlw$���v�T�G�Kn�X�3��� �G�?F� #���1�ʓ�~�~�������v��;���_��[7��~���ƀ��8��D�s	c���ꀬ�vs�(�:�g�V1WC|+ )��N�K_��W����S� �
:���+^�
�w.tDz!����[�x�� �s����LMQP���2YM\9�gK�B惎�Cٲq�!C����w(_�-�%e�"˙�5� �ח+T��5��mZI:�bOm(�C�
�+�D\7�'�%�C5x�~����׼�5~���9���?��#���W�D�p��)/C� �n��<sV?�D�֕�B�˔�q�>�Q����|�����v�;�=�O*����f��Fy�sQdX��E�ab�5��8pa�0.N�Ȅ�� :�s��ҋMS��ՙ�?��d��="�8�5\�h�.��b��>�_zu�s���p����'�p�7i��q�#��{��u� I-1D�T�]R��|v]�7ma�P��2~��H�:�(9�B�am:�]��֬��CC�p_��MS�O	������X���#-�~�z`�`�'b�	C��@�n,|�Z�겘��=QP��Yh��E}���>���6 zX�� PiZ�C���[�a�tZ��:�,�-�d�v4���%�~��*�b���r+����;/v���p[�m���ؐ#���-�'#�J߽��?A��s��\aoV�X�Mb���V6�2Z�ΪR���QIQ�"l Z�%���%���H$`(���P���<S9_��^֠�UJ������S�?($�O������T�q���J�8\`�aa�"�md�cTH�3�9��c40��-���1�?F"�#�R�s�dzYg�]�E�`�ey�pyE"N���yFL�<�P$^Υ"�ӝ��,O��':̾����w��{���<䡎�!�w�����F��|]���{�O�hv�2 ͻ�������$v��{/p"D��q޼es�V׀�qM��RGMP���q	0+��n�T�	�3
���#a��*Ր�:m �v�΢'s�f��݊��y_�D� .G5
ppm4-� ����i��2z��@��#�=n9W�B�G? P̧��x�y�JuL�����Qp����  05����M5�=fVt��N�1gYWߒ��.^��h�����p�gh�R�}���v�#̝���Ĺ�`�@0��s�B9B�؀*����A>�� �?&�C��\����&�Eg��LXƚ�:��!3��z���J⇵��g�C��(�k��:`z��el�D�r��U�����L�?6>�4>�'i����� �Fz'*�|��cQbMB)���	�7�!��Kc���H$b�db�p�r��+�6��qhfp%i�_ w�>�}����U�<�%�t���}��^q�ŕ��N
V�.,��;L�+Wh'�t�,����a�.M̙!��~z�����B�'����
<Xl�F��� ��)\7z9"E����T��ڽ��?b�M��~� B�ǔ��,��2��L���𰢣��.Eōi�I��ԗ0��O�u�K�=�x�8�
���x-W�V�c�b��	Y�=y�&�5c���w���v8X�{L�Hm�o�!���fW��M
�����HװOb���G�h��"�vi�	��V-'L$�#��#��0��*�4S˄��[���[2��燎�x������cj����fn����Q͉ A0 v"�2/�(�y�Ffm�45� X�է37�J}�X�)����> ߵ�|�	��@0N�MhL��qf��� ���2�	�v%$�2���A�ܙ���I[̇ ̐�B�j�ؿß5&��YȖ1��M���戂��q�����Jt@A�ٝ[��e�Ll�S'�7�&����1?�w��)�������и�g��>f�����ɕ~�p�r0Q�囪�G��cUw d��2eCs��Z�t��&���W��*�1X.��rNٛ6i� �������p٫��e�V�Į�r� �6"�#��g��R��ĸtO[�����5=�C��
pc2-�_6.������":�!����l�{r-���n�����t��9���8ޝ	����6�4&^�����xSx)���:�@�����&J���N�hOSC/2��|�k�co�%�Gdg�5��%�h��h10~�e�r�h�X�K
|�N&PC�@!�����H�����Ȅ�P�\�rx�������Y���)��\@m`��,��GwM��tT�ay�U�v�;֕W�F��y�m "x��6ch�RcJڶrx���.�.��"Z��1rfO��[ ��jL0�y&���+�`9��<�h7�@k�d��p{f��.��%䱯�1!}C�p\;�� pFj�0���,�4m�	W��M �;t
�"��j�	�]վ�G;"l;��z"Tֹ9�c;��*B�)����B_G�� �����\�9�9���!�%�W��F>ª�O<f�N{0���5a��&�y\tU��閲[G���?]{�\w	\q����dv��y\�y�e#�'�lK�=m���pvm@n�mh�iQH�YO�8��8+���K��pң��=�� ���l �k2��� ϊ��EYK�ch��M/0��s:r!��˼�T�*���>�A�%7�W��߇�����	�צyE-<�w�ޝ.��W�<�o:�E�Ş�_ ��ۍ�0w��˖�S��ψ�Գ�v)#�sv��4+y�]G._�~獷s��7�g'gf�Q�l�h�li�5#?Z�F��]��g[5�5�x&[�u��\-ad3u<���g���yr_��p��?T,���C���rO��"
�(jZY�t���{���\<Q�)�Bw{A�h1�7���Xd��#y���"H�� )�$l��`k�Ң�-���(�97)����eK˥��3�h���)�V(.F;��~h��P'���w�͂�b����:x�E�0"T�Fl�:t �6�&�ȶ���܄�g��a�C�̮��t��໬IDw�ؙC�[/T�C�&�7��nt��i�W�/ Z��Um��0�I'��y�[�Cl.��q�c�${=ae�_T-�� ��(q��e %��� ����=�F80,�h�ˋ��)-�h� 9�֌/@��XK��h|�0n62�r)�?�I)���+C�q[9^R��Y}�k�e#����g��^�gou��Y��*(��\JÜ:�t�eC��1��f@�4�W� 
���a���eܒ�3˨�H��kFPp�8��P�;�S!���P�,�+�}�o�4g`)���r���*1^ ����n���> @,х��}B[�,�cP��S�M"X�x�B�,}��>�˽ N�4`��u��^�vݼ����pO�7��iS�u�:�tS�
�x�mr��Nڻw�>��8����.�Z�����((A��I� {�;���_sF�kk׭)�y�RJ����'�)4�w�ջ�v�l���)��H�/^���/�Wm,���������W/Q4ٙ�iG�����jmj3��F3�E!�M�OM+��&Mk�4��0ݦ����M�?�z��kVϵbP\WrN}1-Q��9/�ֽ�+JoLc�8BJ���1)VSt�dOg���s�nk����6���������֎�aٝ���W�����-�ց�0e?�_]Ap�o�7����jL?�a�̏b��.�{��p�4^��:��O��4L��G�I����r�5g�bâ�]����
�;k/�=AB3��D.� 5Me��:ch��G*{�J/��c3���/ᦩ�A(j-fֳ�EHu��s��JhBT�=�:��a�n!i�v@ l�ݺ6:tF<��4�S	��u섄ڴ�s�7���w�n�
�! �k��tR���C�1t�c�}`Z���0 /���ON"�V�MW����`�~Kf$��=Ɉ��2� �4P�G�n�EZ|���?���I�.������� \��С0�Y�
&�����&�g �� �2;�a� ?�f�1���8�9���{�o��H�c����0y�q]��\?���id��9y�K'(���_���wf�n�y�d<�ېJb���$���;��,�#X�(&J�16 �F捿�N�Y�-昣/+S���c?��`J=H����b����s��/#�`WiO�DĄ���ql�~��LJ�"c�gn��"A"�G>�>-���V���WX�GAT������5�K`����u(���O^��*S��=��d(}�CU�1P�ʭ�3�� ��b���P���`� lK+�:��&�,���6yy$���w�q{�����ܵ+�ꤞ���|\�Be7f[�ȸtQZ����M���ilxpE�����VLu4��j�X�1���* �ǈ�l��J�6�Ƥ�sOb4db� ?n��-�ss�L���M�qff5�4��f���J�ߥr8����Q<��QC�y��sV��Y�z�����:����,���_Ѧ5��.��W,����]G�{0 ����=�@�������{ � A�OCC{x/���Z�F:=AP��Hbw�k>Z���i��`Ե��������\��oc3k�0��ᅒ��f��j>FCoe���������j(r���	uȽ�{�u"̹2,�wkDD��M��-j�S�t�^$�� *M��w�y�܇������V�<Dh-����O�c.�c$d�_]������^��9U0�)�M�D�Ic`�*����>��4���ۇ{G(�
ظ>�k��� F-`���HX�­�a�9ҝ���J_3��،��γ~z����Nc�ȅ�����`�5�t�L�}���_D����e��ڬ =@¿����2]p��o�D��*�q�@��xc	��c�}g��=i�pAu/ѹdx�+�����!A!mu~J>�0-h��C�S(�:�<��X��p_�F(�\R�N�`6-wF�q݅CF��<�;O�p���>u-�偙��������ј���`�_R!�Q��J�:L�~�`+��Ql�ꜭZ��T֫�TO4�p�_�V���\�A:K	�8�?ֹG�uH7$׹/�\h����n��Zbb� cb���K��2Q*�GJ||�[�)w*�ę���.��g�Z��:N��	����_9�Z �=��|��,�l�]��}@��srtBd_GG�ܧr����=g&pz�)�<� �ʺ��\ϼ�� ���<f��͐]����:�O,Qn)\O@�ǽ�,�kF���}���Z'��Z��o�c�_|�>��"�O�t�aW�vl��4�@w�%,��2D���7�	�hI.:<�Q��� f���صZ�"�Ц(���ף�Ŝ�p�B|����v���w�e��N������f�� ���&��!��̑��7�*�S�T���]ka�VD�z��n�i}֦v���umNXp�Gϱ�nA2O����Q&]���O��1��NLnTF����9G�ՑY�޸���������̦���ۋ�o[f�&$�����ٴ��R��t(:שF�sY�+0�F�Q@Zۤ��H����(�a�W;Ӎ�@1~2:.k"a8.�0�a�X�C�5���}���Na�r���ѷ}r��W\FP%+n�x�[�c�v�v�[)��[��W�^�q��>%�Fk\�z�]D��wiI�Ř#h���� ��M}�J����eZ�K6,����$Kb�
@��u�<ȿ���>���쇜Şy�F��ĭ��x8"K��ui�#�`	`�`3l�
է}z���y�h� �0�c�Hj(�����|�䠿0��7' ��좋�y��Q2�ߑ. "��6�{!���߸Ϙ��p�X���oJ��=�}�Q��R�8~D�d �1F�J�h���N����$�}�ވX�r��(��M���/[�s)G������۷��ؽ�ܶy�A�I����>�6$���թ ����x����H��%K��?��mV�f�VN����Jsrv�E:������z~,�ieIP�X+d����1��ߛ3MaJ4k]l�&bnvttnrj�����Uϑ���Y=6�*������Kc�{��&�=�[�>:x��\�c˶m+{z���t�MԿ����U�����[?��( ��4��!�9����[�Z�o�O�n�6PD��D[���=� ���%?�<���`��o"%=zv�l���ʲ �PH0�諕;�a>�lP������Z�0���h�csy1�
����P�ι��*��Y��ܷ�'�|�$j�a`6�^uY(�b��ϭ� 䗐n]�s��`�O�.�R��>�5����hR��<����f̽A�� ��,�����i�k���s��n�-s�F�)B�c�4�����ǘ3�{��¬��^F��,������r�l��s}@�@���c�(����}�ͬ<�ݕz�������+0)���x�h>Uu�3!�q?�d:���s�8X<�\�+�M() %��v�c���܋��ȿ -�Bg�*��U���*�_}nh�ѕɪ&0H`k�	]�@��Ww��F�4�ݷ#|46_k���d��?�\g<����#p�����ɰP����F\�&*�|U�7@R �n\���c���"���X�ڗ��.�-���2N0�Y0��ʹ�d���pUF�
��u�h?נ,�Sq�ޘ��^vi9�ӜHQ\ߛ��|X �(������;����w�( ��v��Qe�7��nO�t|G�ɛ4�lǝx�˭t)�]�=|�yڨj~(4��Mt<��r�)RlF�.�ы����][6�ݷ�i��hZϵĵL陚��gRB�I����x�֚&�f�:�U�\i3ۦ��o1Q��L��w�A'W	��ix���M�3y�	��
]��3׻l��1%����t� ���Z�w�0�\Gw����n~럽u����*o߱����bݿ�"��u���9�hT7Չ��4U�?/y����7'JF�З����G�"��qg�A>��ߔUD��9�R�")p��
QY��â�wn���+�b�@�*i����L1n����ؑ�B"�v��O���R��0FDaq�v-�?�3,��6x���&��:��BR�Ӂn� 7�lZ�5�t��2PD'�7ax�c�0l, ,89g`����ݧv���0�ܻ��x����ݬ�.=��#!C��r�z̓=c� �H�<����x��y�.��Y�p|� r���r����l�f�[��O���ܗtvi/wV�����iCAfv��ĥ�{��F���p���	8����ȅ+��0����%'CJ�)ݶG���> �ǐ���{]d͚��א'���s��8�Ϯ���ܰ[T�(�P�J��2v�T ��V+���Q��Ԇb|�tP�`z4�Z�#�"
,���5N .�?� �!�$�B�n��Z�Zc��U]P�q�]����'+U�o�����5����Y���Pb��zZ:/����02�>��0"�sa��͑q�0�r��s^!�1�g8�&�m�Z[z� Q��"SN�A3b�FT��4�t� ���޲��b^��
��OP߂kRm��r�-�O��r�
2���)O|�T��(�ץ�1�N���a�t\�Sd�g3�9��}�� v��Ng��3�Ƌ~#�&%zp��k��HC4���)J�g`�&��ظ�5V�]UZԗ�
�z�����Ǟ���֦z��I^ׂ�k����n4��̤��M�O���7�� 6�Zg`�b�0i�]����"jKԢ9�K�jh�ĵ
�=��U��.�@�9m<��z�dwWOc��=���7~t,���G�z�v)L��b�5�'����_�ii���f5Ɖ���t9���ֽ /��7�n4��j��XDxNà����"AZ��u´�A��Ov�z�j-�wo/k���#N9��ɸw("l�έ�̳�p��	r������/�4��W�B߮��42Ƹ�X�i���%J$*�EtF	;�ZK���bZH��ު�\�����l���)|'��}���]��Z�`�� �'��!1Ȅ���h@�o1��++GB�9��^Չ�G0���`mt���ݸ
���E���M�� ��I�"�}�]$����lۈ�act̰�H���U#ѯ����U�(�}?��psoD-!���*A����0Έa�*
�93�zU���.%~rX��^E��ݍ�S�9r��xh����hK����׸bq��D�@����ɸ��$���#I�(pe������d�k%¬��Т�x��,٘� O�h-��.N{��\/0Uu�^&�A ��{l�yf�"�ML�*�@�R
��d���2�#�>� � N�����'��eH�,1v����>E��H@=��`L6�jd���'���$8`*���f2{6ü����L�r1�)���;�|GlƜ��?���7d����?R#�a#Z�y��P��=�y�#��ی~e��T��'����(��L�Ђv�$�=z6'��0?�>���
�ɺթ�3l�p��z�i�"�]wp�U�+��X���ʯ��T�F'٧m71*�t�y�
�t��;�)�b�5��ɤL%�-�z4���MO̖�#x͊��҆���2.W5��1��R韶�ܫ9��)�}�lKSk�p|��X��yP�C�y��e�k��E� ;�#�]�"3c�f����\@�H��c�RT�q��%
`¡l�}mN.��Np�hK���p	̃�
�,�s3�Y�q'��w�_���r�QG����o�cV��=;({�]��ǚof����R��L�����-	��A0�]�$( �T�I����j�s��|�u�T�/"giFt�=TmJ�S0g��c�(']�#��)��ΞϪ�%Ȍ��ܩZBv� N%��� ��YÂ�'�JF����p!dY���@�����[�0#�����$���ƫ0��~l�z��7>F�U�9c-`kw��.�pO��=�q}*J;��q�n0�	��[��t�����C�Wא��4qs�#�O,g�q��!��Pv�T�W��e�ve��Q��8o���U��\h�>� �����qF"B������,p=3��t���6�Y��2����e�gTs!E��'��GG���-�0_�Լf�ý~d���b� �r.x6�{0��#ڐ��|F��vPi ـT�84@0��>�jm�Keu�l2Y�!b>��m�r�hS`���r��~�;���~�Źs�nϣtq�e�Rϻ�
Q�B�X\�f�6;�R.�f3Y�}��$Z�V>���(����Y*��y�:�@����pX��W���wP:�f��1��?0<�~��9]�X��d	`;�Y��Ir-�'h�"���f�������R	0�c�3$X�C��X�����53>�?�|kGkK�X|�T�����?�r�n2�]�Ъ��{��;�Wa����>]�G4{�y�W��3��id�Y�M���e��/W��������׾�\�;��}ʲ�\��]*�x��%���K���͡�����,����DF�pz�����0���+�/�S���a+� `r�ȖcYd#��Zb~�|.$A��7�g�`h��qI�u������LFHi�
,�%Z�~ff!�<5=nj^R?AGd'k�*��v�~j.��i�ÛkVh���/ʲ�<Q+������V�j�|W�J�3p�ErJ��{`���|�`�8b�m�d�Ȯ����"���T��s�qB���P������ɪ
������gq[�}Vn ����ӧ�#l
cn���v���2GM
j�KΛ��J�LH��'vT�^�i�t	�� ,��� #���滙x0�gy��MWZ���vr��L��85A@��q���\Y�H�8>��l}�w"�s0Hb��.8�8��Rk�nK�� (��yfGs�,�\�䍸�����g�O���<��#�$�1�(C�������)�>=Od��(�&J�gZ�y�;�s��5�D�� 7�A��h*�"w� ��_d\S�P��=�
 &oD%2Z��C�q�Pр$`�sS'�tR`~�V�̵�?�,/��y,��� #�2[�W#P !���i�����6#C��<Gw3O6�h��(8e��kWHV���A"����MG������m�*���W��R�WE�[��lF��\��F6��:44aT�
�
(33Ca���`f�pD9�����`���� ���,�hKԧ�D�F߷ؽ%��D��M�^#�j�4<'j�u"jTjH��rB�q;M@�A@��:v�+C�3�s7������ �C�
֊vf����
p�4�}C����eU��@w^���Z;R�5����C�Z��6�Uw��V(�HF�:gT��UU~_�~�ڲ_E_��nh�����?���I�@ ,єF۠
�%��V��S���:��#���V@�h�} �`��1��J�@p�}�Ѵ�#�^��>� b[�6�r��E��7��r����ՠ�K�=/�`��0[�@�v��H��2B�ӦM���n�%=�Pw>�Η:$Y�W2I�+���;.Y����Mmwm6mn�h�8S�����LS�?�7�s83�f����p�n�\K�9qe�s��o�UN�fm�V{~nSh;l��7�,�nf�߰�Q����{��O昂~"=>����b@�(�(o��$�JY'���"�6��Svj�6�s�g|Vc<���-��9�_?M=���h�4kQRГivW�F	w��ŧ�:U/�Uא;�\��O3�n��O� ^1ų,E�� ��������W} �%b�.T����
�d\ݠ��ZyE1I�R�d{�6��{e�:��>@�i�\�`D��ˊc��-'��r�ͅ��X�����~r�r����7�u0�|�����"M�2��8��HC��(���1�ac�lE�~����cXls��龎��n5Y'W�;\��PF�OV'ٝ*V�Ҷ-��Ic�ƕ��}\/K$0p�Tƭ�pfi�"�q�Xԉ#ÐEdQoB�e���p��}��j1ͽ��ۧ�7���q��������A\j?��-�N��?�2��[����z߂i�	lٺ�!��Q�@_�`�����(����ka@r?B�����L� �t��|�J1oӵs5�4�J����c0��c��W���-�E�'�g���"1��<���H7����T��̈́�-T�qnBpK�EC�<�.��K$�H�|��L��������:{f�A�uE};�,׊�& eu��>�t�9��>�ktЛ���!!3����;��c���UXh/st떭���.��Uש���Dc�U���ci��޸�C��Q��U�Ba�N0��P�ճ=FrC2�K�?>AnJ�Dy!�4�"TW���_� 聏��@s-z�%'q"L��w2A��n�L���댙���J(�P���w�-��(2���@X�b�r��%"[/MQ��\t35���ErP�-�݊���]gr���AJD��XT���Ż�LU�٢��źJ����k��b��pa��
� �%��п�{���O9CH�O��}h9��$�^�H�D���<�h�������y�Qdqo����ܹ�~ K���-����>0(�b�Ƌs`4�DaT�!X	X/"~0�yO�fg�7��)�e&��nk���xF��
;�yU�S�g����01��+U�;�9�C$`l|����w7i'����_���d|�\W�Z�{�XJR>�;'�$y���¥O
I)�:t�sNs&Y�dW�7�u�J�M��Ƞ��'�K�{K�"�`�s'��\++�3W���$�LSf*N<�$�1Os�-�U7�`�1J]X �V�[�6	��!�h����\��$�*�/n(߯�a %�(5<Q��N�66G���\��g n�("LٍА�π�d2�����ϙ�����=߽V�7c�w9c;��]�x��;KE��>�Liؖ�y� ZbiF�<�g��'6!�&�#�w�{G�Q�p8Һ�N�u�8���Ǖ����T�C��Q�Q�G�K��_���m���Y��7~����6/���� ��W�`U���Ñi8e��F$Z[/L!��>��Ǹ��H���k���n9�-���.JbE��*�t�_ީň�M�Mc eo�n��7lX�Z=k��v�̳� k2q����ga^4Q$3v�ro�#EN2�F?o7���#�3Z �ó1��� �����v�E�Gj�>L�;`���!ȕ��r׎1d׊�)w�!�U!L��5cH�<�����qs��w3o
;e\9�M:��4�
F�,�@�T��x�u��GD]���	��{�J�����v����Y� 4C�3 �v�H/U���Ũ��Q���煱A�f#�Y:JO��e0�#�0RT
\�("MȰ��w,��U5>�1�6�
�� �>�7�U��?�c�'@Me��F&4APjz	�wj�K�2�']�K(j[�g�z}V�t���yM�$��|���&��ۄ��|&�0�Q��qA8��H�G��O] ��AK���=��މ��꺌	��D�K3��]�^��p��k���2',�w [��;6(�+J���L7X�9E������/��9������˳����v��իW��N=���S�R����9�xDy�k_S��ǖ�|��J�y�}µ��)�7�v�o�ʘ����v�^m��sOt`Xd'����k�1UDf�@���4���ch���s_<�M,F�=С0�A�Vr��� bծ��6���ڨf�^�|/ڤ�����!�uxxB��Ouun�7�̪��f�0���#��L��8(wҖ���	ǝ�]3�iІ���0a��2�-��)��i��\w�,�)`�d�C�)h-Ad��Y>��z���Øu��Zh�m�x�MS�$����0;>/�����!�����i�K?蜸N u��a>����
�:)�9��)����U��]��R���dE��;l@�ݡ�Q,0r�J���T�B��( ���g��޽��h�Z�	���Β|0�(?X�HD{a0ƕP�	$ɩ#P�ѡ?x٠j�$`%�L�Csn3B�`#�k�N�b�uRj�m�Ů��r�۩�NiX�e�n#�u'�7� �Kԝ���b�rӯ���Ξ�&���|N�0��F��Y!�͈�=�BN��Y�q�y@#�E�����@����D�U���	]k��mkF�Yg�4�h���r-�1�FD��� <�����NX�`r���W�缀j�)-���A���xv���W�˦�2 �am���^�(���oh�"zrґ��@5��ɒ��Z��<���F4\��lh�x�6n�hWn�n��|�K_�Ɖ$�0��+��ԓ�)�>����_Y�<?�ڐ�ls^�,o�\`M�2.�aD��\���U�(���i櫊�����En{��]�4cc-���D�1<?��Yd�����R�����1�.<��|8��<P���6�+��d4X�����N�x��Ϊ�׈�����P���"-�9�2X, �S�}��E~��g����bM��1�����ڐ\��a��®��r�	� ��횯
���'��Yޫ��H��L�:/�G�5*+D!Lt�v�]t�Q�h�p��06`alc[�\ 
'مԠ�&q!���E8�1��['�S�H�ƥ�<��g+Zg�<k���2XQJ���|?vOx��0f҂�	��ڔ��/D���Y�7��q 9�+�_wݵ��~�.[ج�PqJXv� kv�w�q�˯�_���j�	���X@p��W�Ez� ��H�Sۓ�FF6�]?v%����6pOb��7���<s���ΕA�mH`�����xS�Eh<7A�|ޞ�R����4�rY����zX:�(�B42�1ܼ0B�9�XZ����F��7��/ܓ���<�!ժ�E��z̨ P���l��L�Y�s+]�#W����bc��s�C_g:�����W��o�Vey�9ڬK�|���eZs������n.?���GM��/+�����*�Wܴ�͜�樲��k�E��sĜ[�k�5���J��ҥ~�����H
ݦMذ�	�&kڬ�Yڊ��{�������c=��=ЮtR�l�vyAw���6�G��J�BR|���QߋE6���"���>�ì<�9�*'�t\y럽OƎL��%&��uʀ���g�񛔊��r@I�f���F
V�Z�Ij9�P��[O�sL����?�]�8�~Ȣ9.��@̋�h�q\�
�05���6-�U��1eOypt	�>@��!3�̤�-�U� v&5�����S������@��<� WU�L{�ݴ~�:�ÕLF�D1�3�(��_�$	/���Ds0T�ci�[!H3`�.3�- ���Ťy`�̶	a����D��F��BS�4P���{�SN-�|�#�\@�h)k֮.6�P��\|���i0R"Cv��1H���bu�o�=�	a�JR�t(;�<��<=	�2�<�I0$	R��ioj[�ա���Sp���Q{ӥh�۹�3E[�MLA2T��t�W��"�/�QE���Q�|U�ZD|����4Z7Ui����i��3S]�m�o@1m��7ne\n��ʄ�[�d�\�J���9���r٥�5Ks�ǘ��H �oc��Зըˬ�\�ṁ��5*���Q�zT������E1�w�G>���g��8��1�)�M��ct�ח�|�[�K..��Y#fH�Y����ISVe��)��O!܌}$���T����6:�18��P��
)�/���p������w/������{`=�!d����f��0v�0*r	9��u%��]���}���K������H��4;uv�,N���w�W^U�Ĺ2��2� '"@i�¸~�r�-���-g�ur9pp�CT3�cK.�I'~l�=����^�Hw������cw��L9�`N�/��<#խ�;�f�G�p�TF$�H�q踒�Bࠍ�٥����� 9��ΓU�'��å��"�Ti�w^�I�1X.�!��kV�I `>iu�� ��0 �n"�"����1��.�RF*"�B�E�asn��V�2c4^��K�>������$ߦ�D�;�\�h����s~c̸w�'�a���`���qS ���_��cv��c���'��Rf������~��V~)D����r�" 9�1��ZU�`]�%�p��U���`ب�΋�ѷ��i�Y?��Z�ψ���չ�wy/s��2`	���[8c��H2�G� ��Z]ɶf	�d���cT����,����A���"����wfm+��g����)�Y����3Y�!ږ�,*����r�E���<�bA������o��Z:�`�g��.R��b4+�:��>F�=:sA}Ja҃҉�~���ѩz]/|��*2�h��'�ɹ�����a��5EO(/~��#���򊗿����Yt\��0���q�	'8���n��e��4� �c�=o�?Z����VE�]q���_���e��3i��̡	Z@��i�]<�ǹA�=꿨΋VEi�� �h0P�����GQ�f�%O�B=�z��i��Qĉ�,ɸB֯ۨ��l��=2P�BZ�ĨM��g!����.���N-g��`Q�se�����M.��AIڪ{c�n�/��{�Nh�)�@z~���Re�Ɖ�����:K��J�����#�� g��5"Q/�?����i���Pu?���u��jakR1�cd*����ݫG\Xfd�kE�+�2�	�5ە�vF@�M�t���0I`c<�q��4���[Ɓ� �I��[9����]�i��/\���!P�M�Mԗ68Z�'&IN�NI��8AD���#�kF��r*�@9J�2�|Q��4������;��A��%�|2��.��o֣�"�*��W+)�Iy�����?�� �e��O/k�V�[o�Q��l߱]�n��a|\�Yms�
x�U��O_r_f�H� �&�T�)=�6i��>���vQ�!��v�7�C�D������h����~ m/���$�R��Ƀ�3Vh���x�(wrG�,:#�H�j~��[G||n�#t�y� m�ڥ����� �́%r�ڭ�����oص=�}B�ʂ���p�X��%��Pb���Sm"o�����,`�Pץ�v��{W^q���A������S9=���^ JPKK5v6*���ٯ�,p�c�=�J���\~�����C4�L�{�ψm:��%��I��lV��K4�>��O����-�~��+_��K��?��ҖY����z �{�E�:�@O��LMj�#uv�> �r������J��).~�]��-�+M��Ӫ;���J���맨A�l�Su�f�iղ#YT��`��Q ��t~������0^	x�w��7N��<�ܡ̬��EZ5��e�\&ZԦH��«�ӊVg��,�nW���ejh����r��.[���TX����fCX�����
����~�9;�Q��� ��ݞ^�?�Od�KA�0u2�T���&��	m�� �&�0yp��>MV`g��Q�WB/�vЂ��S�	���D�������I*3袴��w*�$��Mclw'�E�!-�T>GЬw$�kՂ�ZJ]�)�c*Q1�h���D� ����IQS�\�]��Q�t��b:'F�Q�P��eBQ ���մ�$l L�j�\c��/4#�+3C2��G�&�d�. |���
�?&����9Y��0W\�}e��ڎ�����(�E�D�U��#�в�#����^:U�Nî(E��!ͷ�졿i>G��I��0 �Ax�ߙA�5�Y�$=KRO�{��i�8�L}U�̙�a�@�%���!�+�v^�
�8��Ts��f�/��artg\3�c�N�9DS@�1\���� �#'�$\��+!0/g�gKĬp�{�l�W�4m�UD3���1.��
�d��X~(�
��o�"!�� -�N��ϪU�a��y�� C�U/�~]g�F	@Bl&\��`������V�u��w��{\��[�o�<`t睛ݎ��:��x^�6�c�:ʐua�@��?��_�%�ξ�q�3��H��D��K�lN� ����բx�;4��XݹT�\�����ƕ��6�̦��z�c�l�^���fT�Q3.H���OI,
��@������w�>�GP0?�.5� �w��,L�>����Av�i������;�;et,��ı�-c}��WK�x��]i4��0�.|*�3���2g_���D�j-غVc�EDQ�a�=#�['�0Q�
��@��9g�&��ĝZHDYc��
��e�\*�Č�/:���hV�'��r	s׵<������;P�;v�>�G��4_����@���!�M11��1���8z�� ����H.\�m�jf{��]@��Z%����3���,����T$6���r�KƂ�8?Y��sλʜk%�2��c9GQ}�Q�>�kP�_�t��#�BP�BE1�ލk)KJ�^��-yf1j�u����B/��0��#�ÑV���uּ����c���֧H���)��ӟ���ֈ�Uø9Ÿҧ��f���cT�'�&=��;����I�����m����,]�����q _N����:o��,���d�2.A����3�Z�y��:�s�2Wx���#w"k�W����}���p3F��F��mN̯��r91/�C�ںu���o���.fͱe�Mv����۲e��'�VX��FV�S`o�����������g?�ܥc�D��6	���ֈq�Iަ�����P�%��Lu�Z���cr*�h�ԥ�e����srE�j����63+�t�Ĵv�����Xd��Pk���qF2g/TwO�SC�z��a>47P,���`���$٠F@�2��⸅���f��"F�G��Vj'�e�4�ٶm���ڡ�#.~H�v�֓ஒ�b��S]�����K .���.���0z�J���]��������3�3�?����"�pUw��@������am��`42�p�p�D�.#���A*ꅾ!:y�|�fP�=`90��YD���MF`���,_ ���x��j�0��Y��d|:Čp��)��l^��"�a��\fc�Lک1�R?��Ȱ�����j �=�po'���!HrC��EL�v�s �0~0Im*J��o"�\@-M�$h��y�\ߠ�j���*�9��"��<I�b9�H���e�{�(,��'C��鋨���&���1�莸��?���K.�:7ʙ���k�Pi�s�ŭ�*�
`g6*�;�!����X����ߝ���'�4�eɌy<�S�@Jn\|ߺg\�fq4�̗t�s,�9˼�vtY��6�,Eep$��eɜ�Ṡ=K�*���&�&����q�b���B�\���.���D��>�;���������*aϾ�
|X�qnes�g�6�5-)�;UFc >l������[����|�(�77�8.����Y�i��:�1�S��	m�ȵu��t� ��sIY�98t`�R��-�sJ}�[qh�hW��T_�r�,�~jz`=����W�uGIT�o�ㅕ�H��@t"Qk#�� h!,=@ͽi�o0B7s�8ɞ��~�4���Xt��#]8�Ek%�UT�2�(P�΅h��e���d�V�X%�a�,��]���������0%m������o��~�ca��,��Ļ��棖��.=v�D��sgq�dօ�8F"C � aq���F�v���E!�
� �����L���V8"H0��6���C|����rX���xA_3���v�Ez��q{Tm]�� 3�]w��Ԕ4F�9t]F��s��.��,ӌ���-]nvg���b�*�J[S���8���D��D~ M�j�j��0��Li��VsF}�+��_��U��	)q�ے%��A���=�f�-��7�W� �d�B,��X$�\����P�����\c��%7-&�̃G�P�y�7,���ǚ��ZX�
�/� �|�_Ѿ�}@ ��|�&�L&7C~�v��jɒ}���.�#}��hf��v�7��{�$��h�O��	�U��ʹi+`&#iS�"><��}�KPdrF洳,70���r"D6#0�r+:y�ژu����f���y-�gnV��}���v��G>�b%ʖ�p1�g��
1@��=�v��~�ʿ���?�g����I'���c�W*�ǈ
�H��G���H��m��)�i#�Z��%��̜D�곎)"k��U˺��[�p{"/�~*z`=�a�a�;w�O
��:W�.����?�dq���o']f�+�Ʈ�gk�L�^ AZ�"���uk��O��ʄ��@Yrک��*`P�V�ͬ5�@� ��5b�"2�ňE���v�PqF#*��*�E��L���!���K��'��8\��QM���P`���U������M����){vc\U�[tt9��m�C����'�BAi�9Q5( >G���bQo��2#��WWS�aq��ާU��i&fO��ŵ���^p3�c�!hi�+2��t�"C��������$�CB�>�Qu5���6u����\ �&Z�r��n� Av� ���X�W�(0K�c�8���x0hcƵ���K]-���<��
�e��g�;~�x�"1�p=5�E9�p���-C�~��1g%�ձ�K{`ҍD{x�0��6#z���t�.i}"�LI��p\5�\��}�^�>�3�<�,P0\胂ť�N��3����&��\��E]�X t� �rʬ6�" ��Ͽ���|R����Y���Zh�̮DT!��T�	
��ؽ�`�\D�؆ul��?��C��zV5�hF���.�3Z��Ҩ	���[�~��y���Ψ;�*A��q&(� '��Ji��cܿK�{��n�x�*`c�\_�֬пr (��-�3~QI��կ*�\v��SS�L>T�<����(�LrD�'`ը�kX�B�ވ�c��ٵp�z^Ft?K%֢�ڰ"@�5-]�jtfr�@����w/���]r�T��-�� ���Y���Uy�֟Y�Y�o��̂7�)�д��S��	M>�xI�Zf4W�[�~ǏW{r*���g�A�m�ņ����{`=���|f�MYT��
� �=
o�O^�3�MJsɻ����:�)�F*5!k0��l���qtJ]�x�Hd��"�B�e�G�ƈM�NǢщ���
k�c1����e���!�"�R�#�d��Ι�cM�0<ZP� [N���L0F�2���K<����c9p��`���h�!�(�����5������W�#�\�M�a��y�Aمq����E�+Y�S�@ꬹ��;\����r� ��:�uY�#��53b��D1J ���7 �SQ-�p�&��<�Ŭ����G7l�·Qw�o'�����,tAD�	`�с��l�}�ƍ��E��WJ֗�aE���5R�X8	_��/hς��� A�7�[�Ȃ�5u+Nv��K�]'=�#��~�̒e��E�ʍ*� ��#,�s9�:�b�0'-b�U���rS7M |D����]�k8a�A��2�[l[�P  @ɐ�	WN�����(�f0��i�8�L��ܣ�վ���Z΂6p_��h.td�^|�"���Uq�D�#}�����4��k .r�1��Y��E�zn"�G�Gb�I'�l�\g^u�����a����)�5\W:�BԪ���%�;�Ĉ��RM� ��͹e��}������.')/��&��(���W�^���
�ԫ����R���Ǘ�T/��w��aH��λ�,�����#������	�SoUj�j�q;v�(�(���_#�NmV�}[�P/`ܳ������:[O��;{������˛;�:��`�Eji�v�1��kij�$�eNsxNk���V 3�-s��Tb�	����M�ݏ�� G@�� D���lJSlR�������>����뿲�[��њ8��Eӟ����4)@E������9=�S�ө�����kVi�劌Ea�u�z`ݯ�Z8ؘ�A��b��
�*|��+�`��{,A�}��	p�zj
x/ĮQ�'�����&q�K3���hؕ��c��"����6�v��τ ω'�\��DVZ��֒c2=��H|hL{ئ��&�+�a��Y����p�NWN��|�u̊@�u�rp�(���*�����W�8er!��*��P軴j��pu@��dKs�����t�R�� �Ѹ�����������.2g�óuo� }m��E�w��K�F9���7��_��dwϹ�_x����z��ﳋ���<~�?jv�}��U٠C�j$�f�K���` �B0r��qfgC��#�q��+5jo�r�,�����?�?� P�+5W�b�v ����C��>ùNu� I���+��R~F�p��0&�vSٲm���׳��dy� �N�{��;�� �s��="�l�u��Q㣎9��*�s�]���`�)^:�9�8�}�&
4lA������quz|��LYX����I��F`7mdY6�ӼD��C�����a�m�n�-��M
�1��,��A�=Ǽl�$E�C�2���F*ܖ��(M]�$�ݻ� �����s��\�\Z�a�>p�D\�z~��h�M�s�"�G�[ν]��˵�{$���䖅ɚ׎i3	c����i�֮Y[�R4٫^��r���f�X �$U%���6Z�s��ru�ީ������4���=��G*�gl�4�.��Gu�+�c�Ԏ��]G6�]���ܺjzjNI�ۚU"
tV��g(;J]6�����'F�gD�"S��bd���5+g��h����>�Q������8���ig�qїf�"+��m��r('�{����n�K6��o���s|���`��%7����g���B<�����=���kO��q��)��h�M����G�S���Xf�m��I�f���E&�;�h��Yw�)H]����@Mf�#J
@4ƸG�ݨ/4"��~-<�c����8��^u�D�BtV�_֭]gC�%ѻ]7����8���*�}(�����8�M�\\��X�p�5r�`�dW)�ߗ���J�xFy����ъ0s���.��)��!���M7�����-Ĺ��Eb�H�!�Ɋ��.F{kxԖ��dD��|����+�(�y���6���0,�c�A����Q��N���kVd���\�R&�����w0�>�>I��(w�~���]cD����� �r�-
-W�]p�bV�6co�	��xp~���Gm�a��Z~t�U��`.���$� ��AEf1�  ����_>��f�֯� ���2.v��[�Ns3^��}���s��E^��;�ӌ���:r��&���:ѫ������7�I��G��n��@hㆍ�B���g�
��B"����]C9��ǎ�:d���L|�3��&���3�E�c�s�?�Q�C�P��[��Y~㙿^���'��3�U���ed/�L\���)C��.C�î`��toW\~Iy���]����w���������̜ݠD���3i"Ӏ�O ���)J}�7�"��[�m+���t�m�(��ǟ�T�0�Y�9�!��k���7�5C�l�sK'm����:���.���O�Je>�����.){� ���s(Z`��z�H�m!c�s��bZEkOw�55-iokY��35;95�f���1���l��� �\񘅚_Զ@
?�f�=�����Y.�E ;	�}Nt�z�p�U0������fm�i��V�Gk��ά$	�W�v�ԉg�~��yȐ��_�<p�j���� �0�&��Nv��%2�f��?�u5Z�����P%J����y�����묑�p�X젆{���W䀉�:<�&O�X�4ȏ��,p#2��+���'���$��|��f��ŭ��hHFmH�׺#�Z���P,���hwyAy�;����LYٹ�>~7��S�d�H�oq��� ���4�R��o~�k��^-���T�[���jg]~�[�Z^��ז�?�g�nw<�mP�A�V�C�!D������ �F<JZ��8��  E2EΕ@sx�L���o�zWWw�������,��?+W_s�2%/�B�Ї>ԟ��Iב!�0��1A�=A�Z�'��re<��,�N�`���'�]r%�������s��\�<q��g�"xe}
���c�D�fs�@���x0������p���Y%�H����}�/^��姝rFy�+^Y�h��S@l ��LCM�`.�����z� ��/|W9�|Ԁܒ�����O˿~���ŗ]\���^^�җ���)e��@\��2"��������1F[��`&����Fr7�����gRWn�����<��ǔ��;O�㧛����/?����)�_o��g?����d D�.���[�顇�NųPۑ�B7�3G�VdK�VN8�1�|nڷ��m����"`����/7(�0�[���T���2 G�FBH�k�)�9Aw����t$$�6�80���	7#�0md����;��FH�<���,�|��5kVK�����z��t�4k�7.�q1T-]*'�k�T}P��1ԦO�1����隉���o޶�����O,l���.=�$�?K��sP]jQ+�ӡ�쇤�U�_�!���Z$�-H@���uJhJ)f%�G�꿦q�,�\[�d�@��s�%-�[յ��Uʋ��&1�Mڔ*�������EΌ7ͭP���N�ؠ6�A!�\|ݧXA����� ���Q�U�����L[�����l��W��n6j^EG��W�0�6�����ʿai�\�"�(��:���)�(Hbh�5��x�1�S�u��Ț�Bn����b���t�A�b�]b|?��ϗ�k��S!�'{\yƯ�jy�c��0Y��S2ر	ևQ&)�}�-�_s
��b�Fj�Ҁ(BI�w��]峟�����[F�Mox���*��c�w��Ю��~��_�N1
J���-\��w1,�M���﨤�9�h��\JΆ��~G׃��U��O}�S��`����7O~��o��o����P�0�s��7;Tw�����6n��1�l�w�(ѝ�9I:v��7,��_�:�A�Q����z�<G�v��U�o2`��><��$k����9�*���R3�p}�D���[���1jGy�J9\Z�+��s_��tZ��R~vy�+^%��,3�DQѧ��l�A{QǨW!���! HˬD�	Q7	%J�& �(��/{�����|�|�k_4�x�@ �����	m�/�5�3�� L(�}�.a"@�ƅK<\���nUN�}j�E߇�OpG��QɈ��/��Mo����/}ы�o<��]�d�^%��;�f�V;�ě���E��\	�����v_��.�j<b�._�W�����{�k�����g=�\p�N�@0ޛ����c7��tEE�f���EFޭ���&��Q�ct��ro�_��<C��==�����(�'��D5u�n5kss��ʎ�[�B��|:��qf�z���v�Ye��#$|.eUg9z`E�_�Z˞ܾSh#*�y���F�ygg�Ԟ��wL)#8���ۥY�Җ��`�R����t��^m��8�J����R��n���C��
�*`Ӯu���Z6ϵw�L�(�F��S,LO/���X��4ף��hS_��ζ7u��gm�T���x�C2'�v��_�� ���Et��,����0�Χ9R0FD���}���>�A	|r���?F�J��Q1P��F��2t@�����@`!���U'O�������ߺ��{�x�i�'�F�ta���X���u���r��w8iަ#�*��v[y�{�S�p��	�7�?����'?�I�]Kz�Bʑf앺�8�Ǹ�u~Ƀb,뽭�?ijD���0�P�W��6�����˵W_S���w�?|��G�5������け�#v��=�U��]>v�q��f���1��Q}a��44��	eF�WYk��|����r�i'�����=�}��l�S�����W��`�|5)(޹c���:w�I�9�`�i`�'��:U46D�-����s�9�%/y����֝[�>���O�����	,�r�-e@,X6�����Q�,U@��o${c��@���@қQXV�����ٟ�o~�>�)ǟR^���_{��wV�����}2�u��l�"MX���H��T@@^��WEA�
�Q`���.�{6�d�'�$�������s��$d���/����i�߷�{��<�9�9G �Գn��qt4REc�����5ϛ�= x�!�B�㔜VҏyHB �6lfֵT�<��ԭ��qLz�m۷��o�)��o6v�+_��i�V*,v��a{�8���"�����X?=;Vh�6 nm��B�T|�WB������U�
��mo+�v��!@���b:^���/|���"U��ߝg�Y�d�&m#3�� ����(�}�`.ќ8�e�|�	������2=���?��Ŀ�1_��/��������o��y�p��sŚ5/�{�C��uk���M�'!ǂ����=�ۤB���'��L��ic���T� ��ฺ��:�4=���h�l`S߯\��2SYkv���j�$�j��~��B�BQE���6�Y�\��='��:Ӷڊ3��^�׽���?���Kw'~r|pH&'L:M�s�������$C�$��=�mzJ��(-oa��2}t)�&'���bB����_����$N�Z�ʻL��C�@A�\o6�a�>��Ԉ1���DS�E����m,4��B�U_�ܩ.��-|�9��8�E'�-��N@A����F�~�����[K�����p��X���b"x2+)0(G_��2����1�P�#6}a�:�WT��ب Ԅ�}�R�C�"��{X�������Z�<�L�?>��Ϛ�MZ�y�?����#4]��j��эZ��6�.��b���$����6{-jHN	'ѯ��ze������W_}U���ß�����Oz�Q]��o�-�},�
4�Yt�^�M�@���߭��uFX0��# ��m�7-�����Y����uo|����p��x
Z���������X}�.U��RJ��ߔ�����`l��s{�̨�2mN�<s�����Έl>k١Ř6�~C�z�W�c���\?��O�O�&�(,��~8'�ɣ16�i�TNF*����pČEt��"pxpƷVh�jE������r��,:BcmSذnCx�ަ0���~�Q0 ':��ލ,�����bȰ;�
=o���x�C��ט�P1F�b�,��L�5"p�q�i����~�{����߳=�u�]� ������Q^ &Ԁ����%v5��6��AIF��}P�=����q]O�2�w	;w�1AK���������
�u�c*Z��
�eL]�[1P����9������jD"^�;c0D�X	̭����S2��K=�% �Y���!!���X�
���[��Ă�
'Z�p��&�@<'<���lN?�q	���zV�Q�k����;�����I��WBimhkX�5�84V
�L�h�e(�7X]+18���W麫�D���2�: [a3�p4��ֶ�0Cp�}Eo,��T�i����*`t����z��Aj���P�Dˋ���]����o�@AK4+,�V���� �8�s��|�e!&#��������Ђ�c��]�)�����`�0��!nR�k��#̻��7iW�6;'�`��h1��M'o��b"&���J1�q�&�x�#��C�S��v��	Q�0!����m��N �}Y{x���������`�d�j��{�S��r-�	�
  �	���W�N:�|$�J*�Grue(���7�Q��!�mwtt�w��]���H^��b
eX�'����}�� �<����`���!ާ8C�e���_'�Gv��Z/�y�o�NǴg�>�5����6���֮�HBeez��F��Lw1��i؊�H~:�cO�0^*'K]��}�c�G��V�-��@�bZX  �.�kC�l��Wҧ��O�V�g�LN���Aea-׸<S8�%V$o����#�/0����N�@<��0�ˏ<<F�^�%Y&@-��v?�v�.�[�����/��𪗿2�џ��i�(`��tl?;�����>>I�d@�h�b5c��,-YL���Mp�ҵP�c�ٻ'<�9�o~�,͛�%�M	5��d���_y��^RB����VX`����w6O��x�R��:> ᳔�H��^U4_)��@Mzc�v�1`�9�i	5��!Ȥ�[�f15=����+|�_�_wC��j�|���Zc�E��E��*YA���*��Yi	 �F�QY�:�)���7[� PT-cW���lLo�Cb�j[B��u�is9W�s+<W"�H�om���h��?Z�nU�)����_bd����ҕE��C"��e"h7��l���`���i�����pH5���*6z], !2d���lڸ��/��:�֨h:�CG����[mݟiat��RQT��|Ϳ�vX��nl¹N?�t9�W�g=�Y>�/T+ �c���D�q�
�%=���lI�G��l_��2��Z�'�2G�S�3\pAx�v����`�V%���h�x�'!p��*ɀ*kc���F��[ ��X������&�>7H�0%�8x(���_����H�3 ��.1Գ����m>TҎ���Ђ�:͉����t���b���s��}�mZg�r�SGȣV m�Hzk�i���4��ԥ,5?�	`(^kb��Lꁅ։9F6�O��իW��un����G�-�D��/!�;�}8m2�$
H�n�Rs�J0�,O���/W��6�����p��m��yn\S%�!��5 K�cU�� >���%���3F���@�zC���3��Ʊ9MB�+��2�1�>�g4W�p��`AGSa���(�a�j��Jsg1��J)뎎�d~����ג� g�<�+������{FG%*���8�T:֦M%����IB(�QB�Hy��X�]{wk*S=�6+����lEE�;�}
��ޥU �M#��oL�h(#!���]k
U
5��.�0��o^����[T	�^��AkN\*S2V�����s/8o���XɯG�2������l8ĹI����L�n".R1j��|����<5���.+��E����)ۮQuA,�]E��Vm���[�p�ֱ.�)�4V*d�*ۻC�:��H,����СA�Y�D�<o����G�'����
��;��賐�t�*�-x����S�ozH��zr�i1�hbV���Si��՚0ӣ�
�+�_s�:�U�}Ƶ'�v���R�9Ҙq5��u�pL�� Q����Ub��:OȋN��"6���E$4AX���l��y]PtTI�=,�!��7^] $�&���D�_���ݫ������>��O�hLH3M�li
�[�K����5�Ѧ��	0�S�U��R�;Y�vӦMV����
���1����z�i~��x3�4!�:\�,%���Yx�LӞE���d�5Klj�J�0Ga�`o�3��{D�b��r%�+���c6&M��`0�� +U��_������"2,��*]먞�q=�&��0��ZƖp��C}`�y���Y�(�_�m��Y�К�q��B�eec� J���^d�?�>�yr}��(9n=̖K���O�ح�>�ɮ�Қ12��}��c
�֯2 ��G�,��Y��Vh�8��5���5fn�b霚�V����*%ot:���^r���M��>=۴������T���>[u��������(�7�RY ��%��p�A;I��G��5+$�өoO]O/g��<�I�O��-�,D�O�s�Y����y�G	-U\aHn��v�ko���]�SB�i�
mU�����޿׼
u��x��(��RG^�J�T��bMEi25�����-#�^�ۤ����ᡧ���-��h�?B�I^Y�&��k���0YnҸ$�n�Y����h[�畧aU���<E��}��Ʈ�ƄU+�'m4�����Ru�.��Y��?Q����W��z���z�,;\��hH���w���jO�H�� ��A`�,!s�bw 0ǩ6�!�EV�L�T9٘�9����cQ��"dyHZ���~Y���9}cì։��ԛv_��	��|((�a>�a%�u>���"t34aiuq�m��?�����m�5.������f�ׅ���*L���\�bO����,%g�q0Ry���
YS-QT�ؾ�LiLW�\m�0��{��c-��I�o��ڻ��U��a�{�=& �X��&NN1ǙF����}�{���\e6oTfԘ�s꿥���X�V?S
��m�f�[���٪�D���4�3b\�0.󝂅J+����ˎ�⾱�G�i��c8 �ՎP����5���q��Th���?xP�̈́tB\��[���re��g��e
�K�#��a��笥F������w*kmO�Q�|,%��A�Bb�=*e��Nw^���+Wo
���_+E^i�ej�ºl�R�bq�QezOR�3�a� h����>�|a1ǁC�۲l�Iw�i��;��8����,&���N�N�qn��%p�U�b{NvJ==]��ݠ0ح��jq�*ղs�W=!�Â�%+6OftA ��γ�H�/vH[����VNSG9�u��*v0�B�h�_PL�ea��D����R7�(��O�L�ڸ�T��0F�¸��`_�#$��� �B��b�ttJk�"���:�<�.��!N�D�E���p�������_ �N�<a�s C�jF1V�W�Z��hhRE�n	7�|�;2i|2y8�48��B�{���.H��&��T�>a?>��[����!,�2T���q�F�K�V��< �t
g���`Ȓ�e1�g��f[ݨ�7%˘��\�>i�p�8�z�Z��6U�����LQr@Λ�P�B-���B�dʄ��6������i���_ ,�6,iNY֘��f*�c�b/�f�o��H�ta�3�}b S� ����jx��0��@����;��c�L`��ޝ�k���ya�`�x��t,k>��x[:�g��{��)��8��y�'1��LZsd1�y��z���5UO��m��:�e����Z���	t*�ӔW�3��?��OOz��4��"��)ՠKH� ��2G�,E{8j ��p׸a�ꉍJ'h����.U����p��+�?}�?Þ�]�6�Q��C�5W�j��5�r;��S�m���w�Non���������8�Z`%�DT�ܯ�8}7eU8�yr%W�9�'�\O�N��y�����b�"�E(��'����R{�RT�����k�AZx�G������ک�8(dF��
��g�Lm)�5^PB�8���Ǳ��>&-���>,ɀ�&�8Y,��$87����� 3�]6�Z�j��Tpl`l��Ο�EJ7UU�J[�y���} =
�����k(.��|}�̈� �����&���E�y��X�턔��g		�������cP�� ���غ � �� ����.վq Xb�e�B��\EP�j礔~�����g,�*�Q��|�X��㥦�	�azd% �~��= �ZckU��1�vP�$
��O���`bj~�����yy���,���Ǆy6),g� �̠��6�H�B؀9zqYX���5�盐S�o<'�HxU�����Z��b�3)��@QbL�`"=�b�\�a�#�7@�_�M��[z��S���̰1�P����kO�a/�Y���`����ÊN+�y�� 9p^��J��3mU|��=�浘�5@,F��Zix�u��>��G��j�ڶt�B����	m߼6��٠$�Xd}��
����A7TR�Uޫ����{D)���f�K��![?j`x�KW_n��P��2�!f��ZC���x/�o�u���[�w�7u�[�_�E�XAK5-�4ĳ�,�{*vI��.,f�.��c���X���.�3�"� �`q"L�:�yȪ��:�حӡDb�d-�4,$d�R�Q��Ѥ��)�sBd�>ȓHQ�Gk>�zP �h��筁'���X�V�A3#m4|�
�����u\�.Bl�Z� Mr���!4�^����hw��Km_D��0s���pOW�
-�T�P�L
���xS��	-�� r��p��R��Pd�w��F&��6'�k�Щ�c���9y�S� �rz"qO�z��K��"�lb����.^5�����{������h;�r*�w�
X�H��I��6�\a�O  ��3e��t[�@�݋�e���-��9ՔM��;�s>~oLU �p�Ř*H]� w�"-��6��0cccAz�q�Tp��޳h_�<$�	���XQ�BČ�%�b�*L�����q��92 !��5^��⁉����U�6�y���N��r��A���4R���Щ
	�A�q���=S�A���ФƊ2�nL�kгCr�=�4��o�xX=��q|���Y�M#Ú�B�C�'�R� ^����Eǂ6vT`fh���Oh�j��w�yW8�ÛCI��i+����1S����5>!F����eZ�bX96��*�h��-��@!Xt�m�+Ú�N��W
��BlϘ����R��B���H�@AKm�^-&���a%��1?�1&<�u�t�'��5���O�cL��CN�Ķ��7�&|�+��~;GC� ғU�+�	PЩ��P��@+U1�Qqz�"�+,��\��m��?v�83����. �-b29�D���5�S�K�Q�;:v�d���4=���w�Q�Q���^�	Ǐ;Z�g7�d�=����8Zf�y,���a+@f��^,R�χ&qq�mщ���I7�[�B���>vߑ���5�oK��}��y��7��&6g1h�'c✝��yR[cȘ��Q"(�eH�2�vW[��A��:6 �r��2 �u�0WN���|���SQ���Ƌqdl�����s<����W�M�#� ޏ#U+Uc3��L������yoe)�����9Q�P����
4�ƨ�FU.�_׏��@��n��t\� �\���ay`���J`&�͚��g�y��-3&y8��f�������y�`i�Vx��@��B���)�����;��+�d��٘iz1���e���#���{������.��xm���N�ْhχ����C��F1�e
��Z�\��NZG�drX�yM(4x5g2*}\׌�[O�1s��t��LϠ�V4"�Yh�s���
�I������MX�XNGs�M4�Uv���T��Kf�û8���Z ��%�;}��E�w�I�����T�O� ?���T3��K,P>����ź�k$\v���U,5RFBa�X'�e\)��zD5.Cǭ�-x��j8K�rQ������g�x�p
�p}Ik��O�<R��6��V�>��	���4Lp)�&�[��Sh���5\�!zv�쒓	���u���H�[�5���!��!�P�a�����rᑵ欂e8 N�b61�M@E�0���Y�L�da �*���ļD��Z1,:�o�����&\j�Fکs8���;�.@�l�(�5]�捥�+�Ac�T�29O�lM`�+�;;e9�̱Gc3��D��PQiF%������-��!�gc���³�����C��9�I�	�kd�6Sk�ڹ�Lԗ�����ۋ��Ľ|��Xڈ�f�)~>/>�l��d<\b��f����>~H���y����k�L����C�'�6y�D��J�O!s�.�-I��8v�Ҕچ�4N������͕3�e`�4wKsڠP�Q�w� �|���r�����tK���y����Ѫv=1E��XN�h�fB�F�+��!<%���
ڦ!S��ie���PѬH�R����@AKn ���&d�]��F����+�K���N
(�;��'��6��zBP���m�:wo۶#�t�-V�xÆM�[h�@�e�x��T�bU�%��ߧ�"���]~�(Mr�����ڽzuaB�r��{�Nӄ�Z�y!�MKB��>_c<��zM�`��T�����Cv��A�bIx29m���les���@�ĺz�����!���[@�Wh��"����DƒQL/�e�3^<͏U'ܥ����؝];��p�~���(H�i6��k"�@Hc�ӵh�l=� �Ξ�w�{c����8�t��u��a�)����l�����K9b;��Trމ�I��H�J!90�E �Sf��ya��c�%��J�i� �F���.$9 �Gۦp�}VV@����c���?kH )|EƝe2j�꘣�-��u�35����v���{[���J,��.n{�%��n��ɧ�b�=���O�Y�� ��o� �Tr ۧ��Tj<C���N�iKڌT��P��^��.��k�ǅg��9�߳D�>}��bk27�U}zLZ�	�?Kݻ�p�Ԇ�V�U��:���
1.WH��i*t�f�<cZVu���aeRm��䩭�Ą���gp:�-��V�BU�y�A�9�T�m.��&_���"����D�o'ydX ��%�3�0sr�(i�"SJ��h`�K��/�?�����yO�yh�Ʉ�d1ѫ�����b���J�S�y��y^�M7x4�q���?���Xh�Cc�����@O#a"Տ��ۢAB8pZm�
Uid����mtM�Ky;�6D��Fw�i��8��Y�q ���R��Ս���SB���i4�3�1�U�C=��֠����r�E��:䎒�^��
����Y��2G
��9ǥ��t<��7����|�SB��?���l��{aƔ���U-��ǜ`���ԯʝ���[o.9۽���:Yh3�^�c��6��J)�t&'T�!9H}�F��k���R��f��7�l"�DN���k�9s�~��R`�z5s0��;�j)��MX+���+��9%�ם��� E�DH��D�`i#]��f�lS��������XR0�j���f��ZS[a-W(�ȵ{�x��b �����b�A����� ��Y�����0^�@�?faY�LbMB�]>�;Qǅ�l�s�9�?؁2z��8}�TLP6�c[\I] 
ࢗB�Y��b�[aOke��Q�;�6!��w�czʘ��>)��
��ԉ��6v %B�����)g#d�727gTyZE �1ZZ~c���C�e��<T��t=e}c�̳6+��(p���S������tZ)O_��~o�K2�C���?�[�,2�}\��*5kEG
}����fa{hk�O,���p� h�C&'Y��s��&IG�2���py�X��?�c=�����C| ����Z*���&Y_��[�O-p,v��Y�Z�Ȩ����^��%'�T	���
�J�3V�����Z-6jv*@DL~B�V�̜�ZX�ݠj�̠܍��:1�!����B�.1Z�}��#��4EֿK��t��� �(�6��}^u�uUB���]�s���(�������vE<d�[��<����,��)p,�c��6�)��a�Ү��;��4�d����-�1%�
���s��5@(�Ȇs��S�I(��� ����y��X�ބ�f�,6�e�X�j}�\���Ӛ::L�'C�@��V)]��v�R���!�n\-�-��A0�{���=��3�9�8I��R�?m)|.��plv�8G�[��F�Bx0܋l�9ψL�S lm��,�rR&�EG4A�"�� ~NO8��@6���w�c�%h���Ɣ��զ�N�Wm(�Z��~̇�d�
���3}����SĀ�X��LKgE%��q�Ԑ��z~�<�0�����&"1�)��Н5�as��F!!��R#x1{q�z�3�2�1y0h�>��\��q��L'��8
�y�?B`*�<�k	k׫@�>�bE{�l���kDUC��3��k�)���.��y�Jk��h>w?����z.F���Z:���I���(����
vڦ�;s��Y�m�Ȑ��S����d���'���-��VN��"KZ1��(�Wf��,�S����O��H���Y	SYgi���VT�����"b���G�EbpD��Ic�(k-�c�:蹤�#��7�	�y8�_Rc'a��XM�+^|3��_���'�����ݩe9�˴� �\���:�&��v��<%6�
�y� �D���P;O�P"$��x,����{[ T�gO�Ŵ$�w�'���!N�6�9�h�>�ut|�\x�Ha�8�E;�a7��v��e�%ǏӤT�iY(��R���qL@P�;+G&Z�nL��Ff<���bEa��ϑÇÀD�h˘#n�/��X����Y�]#u^��\��T���#����
S�{r��1��)���4.q,>���_�yĴ`�ʅP�]����=ލ������ d�bj2�(���"*O�!z�U� B ���R��'�Y<�@���S�,L��}��!x���yd��+|m�Zx`�`I9�d�{��Ajݢ�M���p���;��9�9atH�7�*Nb�z/6#TxN��-��9_�b�{�5��bC]/�ؾ\}��<���������t?Sb+��T��C��{(�X���e8��>qn[i6p����2U��V1�C\�l������"΍E��w>���_��Y �����e�ͪ����t,���9�yp�p����?���|2�JZ �����(��z[����Κ�a�������Da�� L�zB�Sa7ճa12��T�l]���q�,z���ݸ�C�[���	�n���K�Z0
�>p2�p8�"CםD��>������)��Hz���iD�]��T��}�_�������*�j�;�_Q��Z
1[ۍ�f6'��i
�Y���r�پ: �2�gi�l��h+�ꌢ��k '��A2U���ݪ��9C�VJ���Z�ZJ���h��+��a���L���c�����k��O���ggb8_bK�%�����&�/6��v)���g؆Q�?�<dU�܉�_<�bsjߛ��q�������!�2�4�&��K�^�#�<��t��	���"|�O�\�c�F�O-I\�7al��&t�:�*zz@E	�l��jz>����f�����,4g� �7��2��'}� ��=&`��R[�poF�s�{���7g� ����'�����w�*��fݪp�m*�I�#5MUx�Fb4]ua�ºzfi��6�_�?[IP?->d� &��7�gA���X`U�ft�I�K����8�悼N�f3Ǳ�=��O^�|�o.�A���=���%�V�Wu_��\ȴb#jYC8#���ÁTjW9<�k,QK�4�v�刔Y���7�q��N3�H�a-��	Q=�s\��N�+����׀ӈp�bW��s�-��M��xT����ض��S8��xB8^�e��x��B_b}��ME��oN =���H��'2L��ς.�ݴ�zD���xD�� �!mwЄ��5���U�uE|ĳ���bz?mF
Ѧ�Ҭ%FG?�g��ɝB�bk @���#��l��N1���38!�����ҽ���1��0��Rkn ������%A��	���iZ���
4 ʱZ��jDI��_Pۇ0���a찏�nG[F����r��=����Ү��j��+  ��?����~M��wc�q��b}R)��A���C��h]�<HvЖj�-����}���4������v���w�zF���+\j� ��F^�M�҂D�R�x�S�����a�$8Osݴ�Uř�+��s��	k�Ú��P�K�]*�A�U����"���B�#�/���V�숊����t~/l��^,��i��z�.�xZ!�.�����}ž����g �x*>"�� h��쏸�f��փ��nYˈ2�	p���,���{�� #�#(YX�ٱAp/�/�({�V��k���1-bc�Y��aR��D8�l�E'!U�E�Ђ�i��Y�'��y���!��qH��4 >@����c�wM�9&�ʹ�Q���bт;��@r2��)�s���S�������<�I{�:4�F[�cw�w�鞽 �����l9�@hA�4q�<? �&�Lwoc����G d 1
dM�p���b>�����U>N��(
Gdl��1�ϓ�!�ᤍH/X;�~1#$a-I;X͝ �����AC��Xd�(Ð�#.w���<~�S�u�-�yikBh� W_����D���c,noS�y���X�L؋�Q�����#a: ��#�Q26����BPr�tN�>~�]�96��i��E&A8@�����]��ەЊdp�K�|MNP���<  �QIDAT����S���;q=p`�l�ݷ��g�{S��Z��D��k�������5Aw٠67�����;���]�����D1��#BK�T���]>L��k��~����>��F�H����L��[NSe�U{�-��RbbyJL��d�M�n��o�_#C�1��z�̍R��� �`�m��-��siZy�>�ZZ�3�_Y�d���փX���z�z�ƞ*�x�-����h~��':�%��?fv��b���0��/���Xf[�%b�#r��ZڲP�*��UW�����a\�[��|��J�E	��
\�;�K�W{r�؉DPV�OM�����(�?�c!�M��0�ʛZ����٥�:)�"F�M��D� -��`��V
��n�r�B��n�������Y&�93�#f��qn�8�Z�=$��އ檌��8@��,~��B�Aڴ��C�EC6O���N.�pR�y�j����J�휓(ݮ����{I"�W�8���W�;D)�ź��rCדBmV����<����#c�J%$@�8de�/4^�NfG��@+D(օ���!��P�s3�/��� ��^�VSd�&�a�8������.��v#��R;3_���� ��B�X	;�դ/r��6H�"5C����z��qc��c@��Y�l�,ܨ�_&\�qM�l���Т���	��;��Xh\��I�gDL)Lt�
`�l��� 6!�K�.�����NaD��k�BJ'�Q��C�:�[6�s�;GÂmUEZ�J�[U�i�1E����Jr*�JK2����6@+�c��e��蔛V*f��Y �]�-�ތJA �5��4�-�;��f�/��� h�cl���ؖ��3u�rl�I�CB�N>��N{L�Ĭw����X�ww <���*��u6�=��MW�֮�V4��?��Jv}�BN���V����$6(�M��$����7c�"��!˚��ݼ3ש5lE��5Pod�p;x?WI����/ӭ\��t�R��yZͯ��Ѝ�Y5^�C�E����4�>�g����2V �{eo��,U^Z+��؀��D`����~F%@V�l�-�8�$�A�P!��Wc@t����������bl�s�{1A��D�I���8l e��H׏�S�Ϝ�ۡ���#��<ܳe��H���V���&��>ll8?����p���3�ź�� �o����Mi�;�is�怋�S�yҌ%͜u����h@���vʘm���.������3N����UșK0cn�q锬J7 V���W�e\ʜ�t���ݴ� @Ș�]��O���"�SK�nѩ��أ^	��r�~�硒򤮕����32Kc�`�V)[��n�:+_���'M��Y(��Bm��A3���=�]ʨ۰~�B�{C��1��Y����è2� ^T��Lu�l��Cp��m�0�f˞��������0tlR�~��e���2l&��kQ��1} ��e��~�ᶅ5:�X\h�3�"Uka[쌀������E��eZ~O�<��֌�k�]��ND��[��Z4O',�S�`��\�pӍ7�Zo��Z��M��,��_�bͭ��k �u�צo��#�a!�F�*Nƅ�/��9�G�<s&i��-ю�z,�ӟo�I�����,�bm�ba,�)h!��n�@��PV���G�G��)��}.�R����M"tc`��|a�iV7{x+�:\��>Q(��A?����9�� d���� |��g��r Y8����7�U��75�8�g��,�ëÜ�@pN�H�9��q�~���C6�sG0c�$�&��YB˄#5]=���H/)��q(��ҢX�F���s�R�;ƒ
�V����@�i���:D��6z��� ���(�%������K`J�o���B�rʤ�{c�q���2��`>U*%�����j�9_	[� ��'d��u���l��`�	����]����`�O�8����Ш�6�� ���`%�� [�P4��0J�4�A���*e�L{)+L(v0���?�;ƛ�^�p�\�R��!c�Rsc�����:�z��G:�5�K�B`K�U���U��9�Ը��ޙ.�D����g�a�,/�j���@v#�xذJ�����ki�`���[������!��z�o�9�@A?���`w�Gm�׌�&�|Bl�A��c�"7�'�;5E����g���g�,{V^��lQ����� �>%Z�U��ږ)�L����H� �3y�������+�x�q����F�H:~w�v��K��S}cq�6�c%P�D�8+q�nF�nD�1u! j�P��"���Uh�?K�2O�aG*��6��NL���VցM�����<�ԑu��������0P�R�q��4 �3�]��1M�<���p{-F��gX ���?s�B!�"�gS+��3���sT��Cu_�����@(}�,��NZ*����*�04��΍��׌5�t�g_"p��&dc�gؗ�U�#4
�R�NF�A�K��ZN��,]��~,�^<�tE�Km³V|1�u�����`�(������З���n�#4N ��W����٫�;K�}�<4�s��K!2�?U}��5�S�i��e�}�LG�G�B��%7�j,;K��2�����Q*�#t�Z)�Y����1��[&1r�Bu�	�Dpl�?E��--9�doH���--�{�l!כZy����h�5�9j���1�k��U�m��P��ιj�
�@kvK�y
�������CG=*��Fj|f�C����S��0�?o�\��]Z+R����y��
�p!��ò�Y�2g<��FW���ߵ8��X�n,�A��<8��J;p���?�i�ҹ�G,lw~,��������p8S��:iE��Agה�6J�N�@͡^�T�U��De��QN�8m	��cD���ءm��"��_zo��S�ARdX,d�\#�!w���P�;i������:�F�XY`�Z��t]Մ��0�U��J�<۝ǝ8H(�ZسYv��:,��$�S"��\o���Y@)
G��l�I��������� �D����v�r4VO�ГbP��;+��D �k`^�%��.�N���c̈́]J+�ؔ[��|<���Z]�U)�ɔ��F�W��zp���o)�1۪l¢.Pij�3l�g��qK���1�H`dʰ7:�d=lF�kf�k�8G����	6�V���F ��Q�)�c�(�1F1�.�0aI��0��s����H
�p��I#Ľ�,�M=�`S���k�{�\����V�-ia|m�fJ�e�����?�{hnn���g�a�V��k�w�
�mٲ%<�1���
�}��{A<�F��8�J��0T�
�ͭ(���¥ R�"g�[�3�3k����������=�ݡIM�a�����+�g�s�`X�fe���������<��P}c+RT�K	 ��C:�dr����0�"V؞)�w���Dz�h�b!V[�";m����-4~�H=��6����-q�y�� �
�}�~i��X=�P�=� ia��8��pG*&�&~�%\_���l'Td�;����v�����;)}k�D�֎҄��Fr$���[Q4�ݺ%����i����ޝ���'T���8|֜���K±,�B�J0s��#�h܀��䜽f!�&��L����.��S,��-A�'��ZX��F"�gfḭ&.�����J�~P���ǰ*��3/�6����.&:&_|u}�Dৌ�����c�#n.���85�4�J���-rL,J��W輴,��/��v�&t��0��s�J�� ��؂6
���>+2*\D��CC���U����������R�Ī>sM�i9dKڜ <Q�,/�Z�;�I�XB��^��u`0:^jN�E�jĪ�q�Cr�5zOE���?�F�b��Π�%�a#��u �E�c�ߺ�j�'���:vT��1;"aJ���(<5*��3A��	�E�?%�P�F	@�XL[�����\���s�0$1m���ha;�/�1X`�*�lP�cY4 9�� 4O���<?z\L���[���v���Թ٠4��5ջ$+�B;��q����y�*K3N�q����@�F�{(�Ƚ�*nj�^c�uo��L��7�>ۣ�����p�S���/�;���#�C�ګ4�4Z�����o�!�ض-\r�B'M�0�~M�w����9�uJ�02@�n�Nئf�"xZ.Y*R�Q��_��������p�:�i� h�#N�<m��P��;M'-�=N�
}��z��G�q�WSN)�\�9P��dd?�l����J�^�0�#M��bѮ��l�L'��%�0�^Rx�=B� ����W-5���s_X��M�������خV��"x,�r���1%��z9&���%���~k/��݂37h����k����d�2�%����;����Y ��G@�'ڒ��� o��uv�ޡ�-4�ԫ�Ƞq�@0�.&鴨�bE�\x�IE%Y1r� کN�����`'l�KYU,�w�_�(ҽ�����] �(�F�0rh���&jt);2'uOh �c�����g+ ���u��gt��'����
�zd�M��5U
}(;�>b3��k|Z����po�um
�H'ҧ��5�Q�l `RN����2hl�u�d�x���0L-�=ٳFA�R��s@)�g�q4��pưڜ��a^��d#8�!U6�5�]�au�t_�H�̙)��
]-�la$�O����y[-䞻��c��a��Uw��������z���'?��p�c��B����K���a�f47p��nR�e�YE�3����fUP�P�xxX̡�dL)��_��	`�p��0^�I�X��z�YB��[:.�@ē���e`�֐�����s",H8p\:�	�|�BJ��:�������駟�ݾ-��8da�;�C_�Æ�kB�f�����2}X}]��w��>@e1V��\�o�>�o�����ϵW��|�������U
L�]'4�6l^jUe�J��<s�
#n7l�g�]��L��, M��z�)�����E�jZ� �G*Х{�>f	c�Tܑ��e�=��j��2�$��J�z��<ОD���e�(��HѴ6X	-�'��~,���a�L�jU��r���^dMw�N��r�H���lh�ĭ�|�C�!�_�1�t��@��P	9K�Q<�
,a�/�8yI������J��{m��P�:>kqoZ��:�[�sm_�,��/�b�-�'2l"�B���Ǚ#J��0�4��=t�D���√����c`����N�3@�}�����ўj�W�^	,��P-c�X&-��9������u�Q�m!L�BY7�;t0Nz�tbӡ�{Ld��ޮ~[a�5�œq�����-Cԁ��gt(?2VSad&u|��͍��;&�0(`�N�YΎ�B��%��d'shC �����tu��n�����2�-��Am�9�k��E�10�D�=��k� a\�8xĘ����N�j��#ǻ����尽�znM���ռ���	mI����nhQ}����}�u⮬�]��(U	��֕X�6����I1���i��ח1W*�  ��hp	ȢAę�/�����1�
�ls�J�h���>r���iYx�s�kl�{�Y�8�֛o
7n�{Nأ��O;=��e/�\~E��G�Z��;wZ�Z���0��")�� v�8���	BM� �E� �ROw��%�_̫V������d@`��z�C�Τ�����ݪ(s���L��S���V{
�J`I�ؖ�����U�t�2��n�N?����jB��{��.{ԣB���Ĭ��5�h|�ll�<�5�]ڗ��v��J,йp�!��{�N�b�"�Ê���5�Ņ
��[o4�����������7�M�P�PW�mf���>)�60x4,�0�Jv"����A�P��C;c�ד��ň�'S�s�����A؄S�S�l��zی������zkk��]��3x������ h�#��S*M*� ��Y����iu&���%�%йq��v ���D��ɗy22��_�����YD�c�"�Z�{^Xl��	Q $���^��A�`ט��p��k��^/}��ڥ���=+,kn	�ݷS�d��;C�~����D�sSr�bW�\k�IV.G���L��Z�r9�Z�1X�~���r�e �����b��W�P��9��|.�Y�z9�>s�k֮7��Z��ش;n�=4�n��8d��7`#X ��=a�}������!sj�C�@ȧ_�cY�L9@�p�T�"�͐�9q� ��a��p��]a@��g�6�_Z�c�n�~[0G�3:��̇��V	l��1��\�#v�c`��/�y 8��Ͽ��O��['��P�0�{F�J���V�����z�5�87�@�m�i2����k`�L:���
g�yv8���6	��۷?|�[�2f�� \z�e� ����ڷo��{��u��E�u�)ï��˃�8&43 ��Ί�0�&h�B*| AXj�j�lܸ�X�Σ��[�V���+��~�/9a͏�;�5�Ҏ]{Cs������B<G�3(=v�[��*5��wBk���燹Ch!��̢�Ȱ@��1Y�ZU�Hk�*�J��V�Bs��H!5l��{��\tX��6Tg^�y�Q"�29��^����� (���=��_ ����>�|�֍ھ��a��ճ��uKT4��(�2@�� ɨ
�b�P&@�F6���G[v`� 3����y�7��C�l/�-���Kuyz�Q���Aa���֬g��9�!�8�£��nиU��3�5b}&�u� �1(;"����0�τ�Q+Ć�͖e�R���bk3�g6���:),��h�� ��#u@�p
�-�-�O��Y ��������0[LC��V2c�g�2�,���F��!4�Xp����%Zt���qR���Hdp���5��)|V1���rv,���\9J���b�ίX"E��#���ж����E���aSxֳ�θo��0��a��[E�2�c�9Ugm�v�0
}N���ؘ�Qe�Q����U|NU����5��iѐ���Ң8A�Ah ��:��a���叺/�^�JZ�M��ۥ]�!���0���8���[o�3hT����u��I�=(m;��?�R�W�[V����^cU�3��u�&BY�6����5�''�3^�c����ȹM[��ik-�����hԅlݺU�`Y��λM\�y�^�,�m�7�:�?��#1���u�Ղ�:.���a�!99&��`��:��
�ӡ����30���E�9.��/�R�FM��2]���r�b
zĜ��|=��~�٦aa�V�6���q\��o�յ6��쐍���}y����cp�IK�ҥ9#�)���½;w�~̯<�Ҿ|�J�>j�A���jc.N:���K�3"�@И5k�.�䒰R��w�����ͷ�e�C؊�9}��v�Ç��l8"�퐀?��"�7����4i�	� 8�ň�ٻ���u�C �F�|Ps��$��n�!��U�����8?JB�5���2�����k�9#pq��C^�\���f.��� �s&02�k���{47~`s�Ea��v�Rg{��}����ٽ�F�ݶ����ф6#e:*w���ԆP�*PI&Yq��p�4Kuu56���L������������G�.t��A���^��&ˤ�?z�Ϙ*6FS#�@/�(����FZ�1���'���8E<K��@��e��$Y��?�5��@��2 �s�̀���\[!TA:A%-�/�O��Y ���O�$���x�2 īA$��,�Ǟ+�L�{ �A�ty@�����SՄ��(��<�k$�C�����������a�������#̕�%D���
����s�Ia]�3�
���6�[�m�j��B�h��Ύ��a	/�8�|���w�1��i��V	����TG�A���F
���D�����g�BA�%²F��19�m�w	���t��"�g�c�(
�>��n��l\���{��9�s�1��o�a,Y5Mqo8�;�u�0A����z��N1D�4�4Ї �H��3�OG1i�t�>���ڑ�����L����ζ�σC dCV=Ԁ�"dw����+׆}���b_Tf��MM]b[z
&íw�c �]��C���B��u�&�(��<hE�(m`)̀ ����lظ>��b��ᬷ)�r�C"��&}8�s����[íw�m��y�i{�ۨ�� �ǝw�i"�U�V���k�B�\cY��Y�ؐ�U�4xͯ��~	x<��QX�0��m>�.�ǥ�u�B�A@�5n�޺�l2�*4� �U�/0dwI�1+pU*���ez�jX ��
����O�~Ŋ�V��@P���a��<x$А��@IG:�E9,V�R�ϙ�n������@bߪ�h��YGŚm�h����%��t��F�%CxL�=(�TS�dL��X���ν��L;�߫����_~�1W��֖Ч�61[Gu�!�X�
���	�ػ���l����(�٭���"��Ex>>�g� �s�گ9ߠ�₋.6�pT��:t��z�}Nj������w&
��1a��ZK�W�Lcݦk]�r�i���s�%��O{��E��r=V���t=�ދ�d�9(�/�S�ke���qڛ�C���bz>�����g[F� ]��{����m-}4��a�Ma'�*-V�-����I.Y<^%�S� E^����bZ�H;���̨��x������V��m}��@�_,�߆��Ц��C,���n��a[\"#�W
�!���_��S�v�=֭�S�PU8��_��R�C9��fD�:3kW]� ]AAuP��̕I��'��,��_-�1��#=á��6l�zn�+�6kml3&e��_��QNF�Q��
?�Z��gF����k�n��.���yv�?��bg�sA�f�s-[*rƥ{�����5�KWQ�p�2|�����D�še��PT�kv9�X�r��1E�3���x�s�㘚B���93eSv�(�s�5�u�ݲ{}x�3�v���OX�v�-�b0��/7�A9��.=˜���L���=���G�K��&��.4}Ǩ�.�,�|Ӎ�5(F�Q�	��u�~݆aL�q�ڵ�
�QШV��Z�P+�F*:E��G=�W��;w)ԣB�
��
v�(<'`�qD r� L��@�L��a�ˠ��bպ�apX��耴-8Sl�?�6 �]����Q1OL��v�ut� �c�f\�k����<e�Be����n^�ѓ	5��� �BF�&P�60��uP�I����U �` �O]͍5������^�98[��Q�z� �v���-l�X�0c����I%psXO�4a\FuM+��5�$� �y*�{׬Xv�Mk�Wi��),x���|-����L��W k����;u�}�b�N]�]�kÖ�N���
3�ܹ�jք\6vR����#�[���\��ZM}u8��L=_�K���!o�!+o�vO,a?ƈ�@2��4��7������y�gP�X����!@���<�ﴍ��F�}��Ko$پ�n��J�-�b��D
�`�K��kB=�� ,JI/�h%#��I^V��e���K�r +����d���8�)��}�c���'�,�`I�_�;�o���]�����+yew�p�V���QQ:' �Bg�X��m@y�@-h� ���p��,a�JEY%VA�= ��uon�!Auv5��e�c1wv��١�ѭ �4*ؘ(�Q��!R�zՑ+q���`h���dVYE	�s�Y���{vW�*iք��7�>�{��fEi�?Zl�J&�܎�k��A�g۽���:���g>M���QN���hPԊM�v��Yao��>���8�so�P��mA�
��
�ᘆ到(�>�����l���"�`��g(y�e�͢l.�A�Y��u�a9�uo��4 �bd*��i�V�S�ʕX��jh��0l,Y|5�0d�Q�yR�Z�Oc��VI܋��n�<B�)[jla��b����@��4�,��u떛&�۶��]�1
�+�k8�a�3c����'A�M�V[+��D�u
gM�v�"m���3o�%�\	a�a4  ��M
Z#X�*� ����PK]�rik�J������_�����-��F �MN��
����55օF����RGH��&���1=�d����)�W�{���y����~�u\@��B�C6?4����Z�	�<����_�П��q@SE��!"̝6�l-�O�.:$ا�Ė�j�o�5�"�Ս��X��p��T]��TM�~M8����ߨ�넴V�z� ����
w���֊+�aE6mۨgz��=��	1˹Wjİ5�铮��4Rht�+��Ƭ�9��iY�|�m�����1��`�i���׹�z��x�6=�6�d�pֱZ��B$�� � +0�l�֋%f^�����j��+�k��vG ��}�����a͖���B禬'^��.׭�Q9MI/DԴ��4W5��U�]�	��L��I����V7K`��Y� �~�F���P6^9��/~�K���U�]���#����	Z�`d�"F�=[�Q6[U���Y�e}��%�r�d�L(�_B�&z,Q�M��Y�I�R�7��Ϙ!��S�b��ۙ���К/|8R�Z�9�q])�U�V!?-^V�_ ����'P�0EA�W;Qj� �����/~�j���(^s���a��i��5�R�N���Z�6¨2���T6,�*�/P�����Ĺ���A�\X?��	�
��M�eF��E�[A����'Mx@@�ki�&��7��bB���ł���Y�&IN}hd�v�V�F�#�u�N!��=��� Ŧ���9Sf��i��ک�>��m,��N�����ڲ����fA׆���9���M�Ӱs�{B��ې B�B;��\v����Dͯ��\d�a�&|���R�� ��WJ��ܱs���+6OʹZ�\�p�"��ׯ�)��p�㺗f�j�n��|V3V�����j��3Ч�V������8&V�g�^����9G�i���Ҁ/��>���{����Wz�54	 H�D���z�ă�֛^}Ku�J���Y<�y�@U]���E5�v��T� SY�`��E�i��J����A��Z� �B���̍m��;�B4M��U��e�j$.�}�����Z�V��~���O���kW��O���x8c�&�Ȇ4Lϵa�ڰR�M�"I��l�� @v\u���Vi,���*�u��5�F����ᱣ�h���=LE���	�h�M� �oVL�%)��Р�?�x����ՑB�s�������=�b�
��y��5�X� Ԛ�����5qwu�t]u5��S���TRA󦦱Ul�6{:�u��T�\�ta��k\�Ț!8Z�^�[�ƒ6(6{����36����\G���v��g��b]�q��Ϣ�%z�_܏e�Ա�s:��z���m�JՔs�|;;�Y>zo��^�a�2MU��r�*��#bK j.(�`x`�i�tw'�g��m�i��%�yq0������L ��e�-
ͱ�.���'TPS�@��Ӡ&�,6u���� �2�B�iRvI��r����!k�X����T�`�hn�U�jG� �Q�'ۤ�M�9Mٝwt�#�#��������'Ѥ��*�!�`P\P�*��8�0 @C�1.`ĊWi�g��,�3T��i��eUZ�u]�1$hDN����V)[H�#2C�D�k;V�� 'ÂM�L�0c�uV��6��s�y٭j�//w@�n�ś���Ε�5Nm%��+�}�{��#�Y���}��^��A?Á����� ����j�j^��ҁu�|P���ѪR"$�g �؄�<$���!2�f4wתHz�={�+�"p'�F��Uh���>���Z<���Zjl���,�0���u$LN�0!��i�FK�E�����H1�U���mPsKU�Ѯ()�Z�!~	XA/�m��C(���
0�ku���0q�	�Jr֑�P܏������|�:�w#b�
z�*cm�.	�3�P�!�^�{wޫ�bT���ׯh����_x�����������}��� 힎I�v��J6ќB�~@�a�&��ö<3#��+Վ���k{��(i�������W���N�  ��DZx � ��!�J�����2�؅�/�jk�Ko��󁭻��t���ʧ<%􉄜��l��xJ�~�JH�V\Y/�'�10�}�2Ϭ_���}������l]@��y5���.�&Ⱦ��q���{^R������]K�=Q{�T��?�c���8T����p��r{ ��?n�o��HhG�+�G�F�w����e�e�=S�\��xI����u��U�
�&XXܭ"6��SoV\[dy��'��%- �0'�����E��Iٶɏ_)�P:ESE����QΛz �R�Z#4J�s"7V,UV�uV�Nj����p��<Te��tl+D'�A�oJ����w�)���r����"�%*�{Wv���� ��XT�kgQ$���d��O���f�P"5�k�{9?NG�Z?���a���#�(ݚ��L$��O�]2�`%��AR��G��<f�J��q@׀�H�`�
 lX�I�B'oB�f���tK3����%���~Z�f��)O�n鼰H�^� p`��(���I�nh�-�u�����wT�r8 �L;�J��?������Ph��<){&+�d��#�
�ɆU�,Ҽ�s���b�	˫T�y38.G���b��R>��%��'���4�G�*��3�e�c��T#�����C�!�N��R�	�CS����z(1D���h4j�_�'=S��l�0��4�$n�@�+�5m�='�5���jn� 1o�^����qB��i\'Z<&��I1����m>' W�y �̧?-�ᖻC�j����u�ݖ��K]�k���c�N��j���� �ֽ���?�� ��j�6#T'W�����zF��}�z�/��n��blm��m��
mP�H���p��������~�-��}��![�ɥ�O1G>;55jʣ�r_W���bw4����Ш�$���!��K�XW�֮ߪ5CϦ�%
��>Q��8�M<�܄	%�LJ;	#&��ǵ����JI�C4�lMæ��Xu��R��V�	�]��֎n�.!��-u�@���	;�
�J�"��bI���^�OG��90>2�qΦU?ش��v���%R`rQI��R�0Y�{���M_��ܾYq�6Ux.�]����/��ɟ�"�e��"b�����Y8��[t��P�E%ڝs�T1�!ЊH����P�X+I���Cr�X\��lrH�q��!���ӄ�X�tl2�X��#��1�yL�"��U�J���Y��W�mi�qܞE�NSM� Nfwk��C�2/�F2��- h����G�HX
�E�Q�d;J9D�t�~��$���B�7YNUrB47-*��,�b��NDǮQ=�)�!�v��$~ެ̰�sq�>MM����N r�.�$A�Ϝ*@�XE�ESQ����K��
�9��z�{�w�)�:W��
z��.���µ���v`�I�19	 ֐�8��u�J9E�T��"�;TPAGR���<+��������0����7���z1d��l�սh�Z�B$��'��1):�J�Ep��
͐�gnIcf�`�d�i
jR�ܗ��F�P=lR2�q.�~C����8�3ij�=�����E�悾����� ,�����o0�:���<��݉,l ˓��ނ��M`�*Y뺭O��kա*d�
9�����n���w@�Ds	�Zk�}˄�g�_��5��CK��0��G�cD gR�B�#z_sKUhY�Y��B��W��ZB&�F�&��V��a/���J�̭cS��J	��xm� u<o,+hgh�f�|�ќAW�f�N�ذ^�v�6DX�&��q*��MU�*��-4��ڍ�	(���g,uz(�)FsF��t1����=�7�7�Ċ��k�l{h����2�jb�YI7��_�K���f�M~�탘�T�׼� h�>��s-q��H-1��Es�,�z��mV@�j�XW(U��ÃS?loj���s�n���>��o\�姉�������ǿ���m;�ٴ|͕e5Z��L �E�(y��iaqA�@t.�RMML���"@Z���vr�_�>;s-,4�{f�0Y���J-rr���ɍ[�i-A���-H�2����)�c�v��+~�K�y�`q�9�ݡ�l�53���f��U�f��Dt^Bl�׊8j�c���9���*cD�$�K�[(H�RݏhM�A=kH��^��҉t��#twxի^^������S��E����ƵXO�!6����ƨScV�=:�.:��g�u��0+S�0�����{��������D�K���Kd�XA(�p���Ӻ� b����e`K��Å���t�ւ6
hr�o�ճ��U��9�Њ�6+,R-�S �Ze�ؘV�8%�K'R�g��)Cԫ��ӷl
�}�U��k�PTqL!۱���w��бgWh_}��-6T�G�ޥ�K�X*����@۴'_�,\��a佧ަ���85i@h�`U��(Qv��h�&���7�ڛ������;?�jOBr���E�;����M�F�C{�RQ_el�lEI�j~r݄�d<J
4J�Bo��PDhXl�ب��lP���$��K�Q�����5�=�Lْ#W*oO����y�y�H��F���	�qғ�8���u��H�
0ʔ#���S�1���NN�R��Q!WD�*�sT	
Uu*� ����I�I�C������3I ��}C��������F'�͖
C*D��m8�|�R؂��f3�Q��PU�jE�oC�u�ze�q٫B���m%�U�1)�6miVv���e S=�T����"K��	�I$nl����MIC{4'������HF�%�V	 �ia��Ȅ���c ��S��:i�3�"mh}��#�-q���U�(���`B=�fT�g�E��x`����sc�u�c/��Ӯ|��_=����>�s=岭���c������W��cfr��u-�[��F�@� � vs �a����@��M��M�^DΆ;;����yfi�����C�����)ձ�-�d�@����xUW��3����(�L���0��݇�!4��ò\�?v�4�� ��1���$f�EP�2\�8�Tk��(t�29*~��w�$�	NNN^[?�`���X(��P�A�����B�����w�����Rײ��*Ԗi���n��J��,0l�n�*o�H�M��p�%熿����xs<�����W�/}ɳ�{�����w�9F�/z��Z]�j�()U8B砇�Ha�RR���5�]��%͇X�:	b�vT��������+X���H���K� �H���{��<�R�ݴ����r�aHN��da`% Δ셃�ƦgT��3������g^&��nQ�ot*�/_��+��e��-���b�z��;L�������e�H�=@�FNw��`-�A��8�R�$(�ac��$�U+���k�B�:=+�1+A�c�?=<����L+ž��o�j��� a@���q��Yh6:кh��&�JJE*��{ի҆�zN�Ū���U��V�a�Rl9��%b�F��Ј�B�z1A%
oRJ ���M�YԼ������.����A��x�l%�����%�O}��#�_�R4z�~i��`6��o��+M���i�
�XSY' 0��-S ߦ����-�P.�1�9�f�@O�0jU��,�8e{�T��\- 3(���Bx�����J������|���ZD=bY9����!�]�9��ӞeD�s
��
4�c�
E[�ѓO��4�c�=U3S���JU̚J���3�:F���pkQESc���PD�?=�\���l&YGK�U�R6�I�4�+Y~=r,�A���+�*�BHG����;�ƪ
�3e#�{�?���=�?~�O����<�����/�����>���V��u����qcqiy�АsJ�@(�"�>�yr�qk]�&���܃|P�v(eCXj�I̯'�y�#�9�BVR���N�[�$��ΒF	0d9f,���̑�?޵�K�������[~�Μv'���C v����5c�p,�
�}���6\G�"E�S�e��]��ء��w�#���O�ݥ�|�$_��ځOJ�FOW��� �i�(t�0��s�>K������3���
&�ʲ�	}��xCx��n��a�V}�j��U��M4l �Ke�v�
5��t�eM�+�k|M���u�BG3�N��&��rD
��\5u-v�8hvχ:K�T���ׇo]��p�_�u��n�fk�4%�4G(��x!Ҧn�2�LY�d �}��_�w�T ת�������7�ax�K^������v�Cb����e��)ۨI���Q#6�D�nlb0tv�W�N8C�)1#ԁjV`���!����0�K�/XIfϘ޻R)��׭Rqʃ�����^���W?W"p�ilJ��T�`ɍf��w��$"G�"�3�kc�
շY	b�W0!��ݡ]"�J��L���1?}mh����J��B �q�́tib����Ⱶ7�Vb{䔩��Nh�[!e���J6+誘�0qbfaa���my8,�${�H�^��/���H�ޞ"1.</��-�T�[��9���`=�R�S�Y��=b?�:P,ۗY�:K���ժk׈)�D,=��,�^� ��3�%J�� <�P�-7�d�A����V�}g�*�K@��U��:ZH[�3�?������#���^1�%#��h�l}���!���`�Mճ"F{��۵W{;�n�����<}Ǻ�+ƚ�jg
�`j�thd��Б�u��x륷o������Zժk��Îl�h����tI%V���W���_dd���#��A�&�G�@���Ukg��Xul�o�+�� @K=<�{�+~�����'�����ӷ�{A�J��i>�ř�rP�-�ژU�<���@�B��5[}g��8@��~9SC/�Ң�o�Zp�ny�ߊ�R|ֲ�&��6��9�nN������S<�Bv[��On� =���뷮�1��Q��l,�� �5&@h�� ��rml�7���S{���p��������K_������:>p4��e/��_���Kj���#ݾM��cd���n}T�I�X�(�N�bAtlٻC�f�s���tw�{�zo���}��t"�{�S���,5�����M�W�P�ޘ�12�{�(�?�q�j��L��.9�^9��pM���k���5��}t��{0|���+ܽ�#,_����;���y�+�o>�2}>�׮T�Φ����-pTר�r�%���O�BS�:wk�,�I@c�t�e��F�~�����o}�{��/YX�^[����s^x�ܧ����`'%����d���#*�)=�e�����Fɡ�Aŉ�.k7�v�U���K�^�r�j�	� ,i\���õ?�>l<�B�v�?��Ԧ���<�4�yv��*2��wy[m�����z1����{Ͻ�н��j[�\�Ju�UȞK1��6�}�c�)H�ݩv���K$EQ��|\�d�K-�FFƄ\��&�� Lw�ҟ������ĳ�۰ hD�ٳC+p3��	�W� e�)L*�/@SZ�vb&���bCS�1%oH�!BD��Ӂ�#A�-.�(��Q���E[�9�?�i@��2z�}?��@{C��6���Ѓ�6ǀ���y(a!HA�bk��ƈs�����Ԩi�*�R���\��ª�ƙ�#���ɡk���K>w��gw\v�9��j��W�x����7�������O߹wە�U�6����3M"IK6��^���hc���=�Uy�A������*rTZB`RMcU��*�`��o<�O8��%{��^�����������γ���G&��I��CFTK�ɢ9Xd-ƄOLc�e���2?L0��ϩ����=h �H��j-�P�T�M7�EU��E d`v�H����r�A�[=��x��p �� ���4u�jت�b�l
�pa�қ����
+�|��v�j�g�Q��y������^�!�\�.�;��r寊��	��?K�'o�hz�D�[Z7BNBK��������S.]�/�5M�>��)�Q���}�#����=?<�I��=đ�E1�hj��o5rd�x���o<���;W�(�q��_�!\����Z�p��ݱ-\pچ��J�^�7��p��#�S�F+��څ��g5G�f�^���A���w�X[x�h)LDd��l��غ�#���Ĝ�fmKh^��å}��d	a�F�O�{��Úֲ��n	o矉u��9�{�bx���+��u_h���)W�⎳r�����Ӟ���<Ӵ&�r2���uN�K�s��yW(]%݇2�i!����רΕ����CaŦ5�}o}ChR�>�@���p������a�u�	�^���7�!�s������GՒcm�R] �^�ꗨ��y�O��Ca�ڻ��٤4n�kjL� 9!_!@sF�����`�I �}h�56�,%c,)��K0�*(��ΨH`��ܻ�Sn��s5�T�.��W�iVɊ�4}b+��dJ�A2���Ђ�����ssT*�E�-�+A��K�ä���d�lލ ͮ���vRT���2�f2���:JC�ź⏰}��<�������t^��h=�ةJBj���P�6�?�v|a������v~�U/~�?�����`���u�����#���S�zǵ7������W��h�|�-@+�r�K�Jg���DN�>����B[ ���qs��b��)Lq�*��F���wΖ=�[�p��PNy�i�&?���^�����_Zװ^���5�N�e�K�-H,Ld���n9�](,p�U��C��ve�ŀ�;`�'<B�2(~���"�P�|�˜��`9v��G>��9��O1c�5���O�\�:͋,�.[4�BH�L:1i��'禦�hg��R8��&��Ii3�شY᫆�Û�rL�r�ii�� "�ٰ�4���fhZ;��=�B���%DĈ�gX�R9���_?��bk�@�-�0+A���m��a�G�Z�,�v������?+���M��кБ^a�����ó�����B��~��jG��w^>���T�G�f��?��й�@����
e5�z4��*�������+_	{o�!|���~���7��]a�ڍ��mM�PhQ zv��E�VC$_, �c,�V��B�����g�|�\}G����n�>��+_��/ޯ��2��,���3����?{G�O��^���
{��1`R&�̊u��WVK]cآjҽ݃�O�����fU��6/��������uo�sc�fH>��&��pX�U03T�T���H��W���rI���g�^�����w�W���I�t(��Ya8��"]oB]2:���V6oj�X�j��@����Ⱦ�&Ҥ�Y�M���#q��-�䖨@v�\�	���l��704h�J4?a��q	ݩ9T$FnRmHJ�a7;�J�G�
<jnQ��Q�7��A����S�1m�B�ZS��u�QE�z�}U)HE	��u��!�R�B���e �A�?�@#��A5%��U��R�r+H�͖aR�Չ�!����r�K� ��ځ�/��/��<���m������877!�^}���s��}۾��?�����W��P�M�{��+��u���_�F��z�LmE啥��zq>�\�j��@�h�z�:)�Y0��e���8��R1�.�׈�i�3G7l�r륗�G���z�c/���?��������u��P�ش:�4�r��Ce�^���T�5jk�CK��(؊d�%"4����x�hPh�rJ�؉l��C��y�9L��(������8�]������d1��Rp�5�MƋ�[�U)@��QW'7�jv(ح�e҆)������r2�^���4_xv���1|�s_
��5-mZ����~�V���C�Eg����Ec@�Hv�@�R�9��d;��ü�j�N��fF���i�bYښ�;��D@��h/.U��ȑ��O^��v5�<+\{��f�"��Ғ�>��S�WJ[���I�&&��k��?5%��]�+��T)YBmX�a�|V06�H��ck��a+|é5*xX"',�	�'����c.`����]�#1C�}��-E!�߽K镵���RS�4O��ϐ�'V�t�Y/�K��"8��S���@'�R���v�]�t15n����v����F8c��p� ]�J�ֈ��߹��T���������7���sT�5�?��7Æ5��%/}Q8����WL���px�!��t?ý�]W�.���S4@pB C�X) 6Ť�+�f��5]��U �u���,$jb�N��`d{�����������������	-��հB-?��j_x�c��s~��7��$گ��y�L?��o�Z�4�:������e�O��X����Wÿ}�;��M��J��:�ڀ8Q���ރ0�<Idt����:) co+H����R���=�&�R���x|�a���!CO�C�V�-ٚa��jp;7>|d�}7��ן�/K@i)Y�Z7u�w������~���i�RQg���峉cSS\4��ʰ����z�X ��%�Xq1ץ�5�%T_�ҎQm��W�Yu`Yk��{ʏ�7U�}�_���o���TQV(�)�<��11���G1�^��91��a�J/4z���!=X?ö�H{u^���([�f���\�cD7�H_����lV��W���#s��}�b��!}OE��(ѝ�BI ��_֗�����FJ-� �5,��Mq���}�I�AS�d@!���u�y�I��Y�Il����%�zZq��n�M� ��S�� ��E��0�.�Nm8��aSb�p*M �V��febV�D�pX;2��VP�D_��T��	���� �`Ũ�\����e:����B���H�oQ-�Q�
��+h+ֲ��M�X9s��,lC�i;�h��; �c��E�d"L��I2�>_5a�}/1.x29D��*�?e�����~�]n��Z���?��M1�%��mo���4f��*�z�����Z�P�դ��
�'i�z�=���}���&�J�2��N�uP��uj�Ю�k�u�Pxޯ>9����V�RƔ�A��3�S��x��qr:vk��m�d��jt=:K�M��@�D�d�Uڒ@���(��H�6�g"+B˦����)�<)��WTo����/{�uJKT�l����ܾM�������Nx��_�'K�Q��^��g��3GGC������hoy�o�']~a8���孍�O�������*,[���Ԍi�'toT����jn[Ɯ�uϱ��^�\�MKD;���<E�����+UpN�:�ȴ�_�Y����P��H-;�$P��Ա}����e�7^��������	�4��l;�w���|}wg�	�וh@�z\戴iM��ދ��tCsC��ʯG�2Z�PKkR�Ƿ0�o&� M��TZ<�m~Nu��5#���t�LU5.� <Q��=�-:D|��ҮN�4&����,	��D�������UY��.O
9���M5"��Z[$��ϧ�M)�FF������a�i�3�@|Y��ź�������:/���*1?v��~c��-&�,���c��Bנ�'�)�R�n\Up�
�Y��@yJ��
iy�%P%��J�E�[Wj2ߨ�LM�&�AT�nN��*9��/�<������β�.P���~�$�8{U���������:E��:z�'\t�i��xr���?�.���]7�RCQe")ck@,@��#껥�Sa��}aBmZOo
=�#�y��VZsuX�j�	iv(<�b�����!�0ƢT�kt����͊�������0pxO�~O�j��+p�c�3�x}��KU"�����sW]$2�&n���oSH�����o�|�+_����1��*e�U��BgBJ�D�N��
��ѥ��-ר�K��\�
~LvV=�9k�Fh�E��9፯xv(��K_�O�lԉ��5�ۤ{W����zj���=�r ���<)��T%cx9��N`uN�ŀ�u�91�cbR���y���۸Vۙ 0�*�N�P��(ܥ��9)���~�������d�}��Xs�"<�O�G;��V�ii g��p-/RE,U��e����j�Eg�_��p�~'���.�������/}~��u�B�X��7u���a��A�c�&�ia��,���,]�&���5��� ^܊��w�	qK�}Z�i�&�زT�Hr��@0h5U�Q�9~��_���Z��33~��Yk�>��������ǏN��Ըk�@aXm&um�V.?��+.:��Z�i��e���8�J#(U�E�]ԸjXXk	=�!��]��c�V�]�lY���љr�j��C���8$j
Y�eb���0:z�0�ؙ��E���%�U#g�y�f��v�Ľ�j�PbV
u��3�@
k��=�x��2Y6��f��˳P]�t�����ؖi���b}RA'_�-��E��m^��b *-OKS2��p\N����XTH�J���P�Be�P`pF5Z&�f�Ճ���s�*9�������.����W�vز�p��'�[�.\q�����P+��yn��I�R-�9��Ë^��p�Ĺ4�,x��g>��Y!���J��]L�\/����u�>d!��=����+����S�|�z2u�.v�j�9L���fi�:�W������<=��տ�ᣟEu�T�*�}9��B�2sEL��g��۴L�������F�Gì�R[����/�M��� �&����Z��OSGt�G�~�O�nTO29ezDU�v�W׹=��c��5k��K?�9O�T}��U��oڨ"��l:<�O]~I��ݲߐ�q�T� Z"�u֨��a�lQ;	F���U���O����7�Is}<��^����	�x�3��V�Ԥu��c�X;'�w�Yᆛn4�UӠZ:�}TF�Buu���I�D��i���U#���c�i��<&;6r8[�,��hH8���j��>$�3�;���/c������"����(|�k���P֊����@�\
�JCF����>��de:mE�Q���d��^ce�V-%�@f>Br�� ����db		��7�m��&�|N��"��֍91S0@V�ܞcv;�A�n]dU�았c��2sMdYJI֖�p���G/:s�w�ҋ=���c.;��w~���޽��%�EEm4��� ��fKssg}]Aij��H�@AKq��:�׆ʦ�*k�gkj�TA��/�^__=��ֺ�P�a:V9|���+�zm��� ��r_��:�	J��I;i����fd^Y�j��H��qzIb�x2��-zY8 ���\L�1L��"ĂZX/�q��9i,���߳xG�X� ��¥6L��3Rd��RS�0D�e�z�����/�~�^1
5U�{���a���hWh@�jU�E���\EMK�~������-��ȩ�y�
��1_�}�=�{w�{�_�W�.�<<�����G���uk%�}ax���rd�O������?�����������i��i���֨�29���%�	�� �t�}��36�7���w�o�0!�J�ݏ)3��r��ן�k�z�w�R��kTQ m�M�cs���������~�	Լ��oox�)%ۦz���o}�����Mi��¯��s����*�o\6m����o}o���[�*�*}���5/��ҹ%hWqD�ղ�5����#��'�#v+�uŪ��'>�I9e��+<R#v�4R��G�7���p�B<o{���.:;4()�C���}%|�_ ��(��������+@��p�c.�"��fX�b�U�P=�Ç�����û�����������f��w�&Ӕ£z����JV�#Z}�F����ׁC���j�F�11B	�������R��Gm�:�K�\����|�����ד��87\#���g_iMc�}����];Á��l�B�z�+��c����k�K+�*��z���$Q���дl��Fa1<�^�o�.zؘ�獴���@&(��F�'W�¨ .�iJ���H&��f���6��6��
���%�?�v�*��ѳ�I�qb|lv���г��巜���a%������?{Ƕ=�zj
�mi�g~b|�\eH�ͯG�2Z���ӍfbJ[.�?* 6Ewg�?�/d-ZY��4='�ش�m��T��vw�ۍq�А�aZh�u�R��X @I� Z�s�vr���s����i�`vX�-x�ύY%�>�=\P��q��t<�Sd��n�ɝ6?�5�=c%~o���YϺ�B�rk�x���FAԺ�d��@CtM��M�x��_��K8[���(�Bw��51���v�h�CGyRn�!T������{{�����B*^XQg���9	W5�^r�.�,|��__���TO�'�/[.�"��z�5��f�@�ֳΑ�����7��@E�ո����O�2��/��Cuk���g�-|���}�ƥFm�����װҬ��()����f��C�?a��K���/;��� �؃��1�
+��j��榛n�ÁЮ����ub+����w�{��^ۤ�}(|�[����&ց�-b�zU�X B�c۶{�U�4�z�/�N[;������תN�5WY��J�`j��À����WT{K��	��v�����ưf��[K�^�a��Χ;l�z���(V���e�[n�5����^��ɑ�*��ad�/���1<U֟y^��W��z��ޫ_.{Dz9Mx�<����QG�X��	w�)�TL�OM�A��A[�A�Rޟ�7�ĳ+?�,,�9�~����\�r;�3��_$|�o	�y�;�Y�~t���[��Q6؜�	��7����>�#ij���G�}����\����*��y_�k������� �Z�*����Z*�@;ڕ��xf�g}�.R���H� �����Ș/��� �_�|��A�H��^�O�o���Os�z�����g�����i텖����usϷ����#`�($������=(�7�i� h�#^_Y6�P]=֧�j�4����?;6��C4�B��K`�|dx����a�����j�5��,K �̞��)���Śth-T�}�Α�d8�q�\�`� cb`}e�(�u<��[w�R�?�;��$/ X�^��7�C�p�m�*��Oz��X?C�nBl�?�]-�ֳ��S�J�+`��&g	E�-��fw��h�-�L�/-9*��D�U��$Ǒ�_���:
v�����W8�P۴v���[׋��Bp#�1O��TEW�;]Yd�]3����&�+U��5�\�i�P��ມu���u��LZ�~U��g>Y����W]���:.��:��]�*�)LԤ�mZ��� ���kC��c�����H h(	4 �%�2��q�{��Δ���c��l��F���.�ތ���OA6Y�v��:��ڿ?��O>��9�P�@�r����YL�@�!������8�f;e�0-ب�Ya��Ȝ�T��C�����}Bb�~b���J�g+ugH@\������9��Q�#TӤ��B{:�*��CJ��;��3'�9!���	4�gk�ig���������m�jR�����������ܘ�}��5�	���i.��>�*Ǥ��0��I��'�M����\`K��z�)�b"h�2.�U�bm����b�fҥ�{���~�b{���5�ݰ�ĭ�Y��|�[
�Մ���{�%gn�����}�>e�	$��	�o:csht�
�\mz
'��5F3��ఴ@�J��Hi�8BN�a�_�!a_�"��6ր��=v|��+�'B�V�Й^��jc3�(V�.Ku�`KƫѵL�ό�jm�XV���"Pnjh����?:��hlvV�
���R"�o��U�w���89�#�j��/�2Z��{�����]�����OL��JX"fw��>�ǎuu������*�7B��19��ʡ��f%r��j��,
���*U�&������B��y����|�Co���K���Vq���L�$�0k�
�-�u݇W��wa2�����r��?^�� �|wy@�tG4t�b�u\�����3�SU��2`9:w�����Mz9��)P����b9�֊P�{FbVB��Q��ڵk����b��u�	��Q����я	�VA�M�k�-�	��7�7ܭ�����7�R�z5-j�9-�M�&^���_�e�!Ԫ���Aiu����0�~i?2)@7��u�)lԶA�a��l=���2S��{z-�R�h���S�mB�U�]��B= ���IP�]&��q���A�]��E��� p�a�:����B741%ӬG"�Ze�+���5b��S�eU�VH7T+�U�̪�e�Y�������F]v�槴�5T�h�
�]r�a��X�\v��Om����@Wݭ���-��ebT�x 
�~d(��e�~�A�"x0?��Ig���-m��B�5�},��W����!�z���[nW�_}x�^~빏����^��pݏo��f�AuuJ�Ƶ�ĭ��Wx�߿6|�K熧]����k���G��_c����pDU�ר��<������0����0���b�0C44�`:�ɂ���d���'2�_f�4�b���9�$���ª�MP�G���*+����Rgmъb�j-��*��..���d�b=Uך�����q���;���?_� h��1�4������̩u3�h��f�;g�O�`�4��%����������-k�X�)pg�yZ_�p��5|R�Ҥ���#���"���3I��=�~��,�'���v1�J:��?�Z#'��������I/�O6�e�&�FJ;M��=��`�F0�X"w�)��	 �杄	[_D�����|X��!��<�rR���c�G ��bu(�V.&�pwo���l}��tPՋ��qf觞���5ᴆ�IZ�T���%�ՙ���������Ђq,�c?,��m��L���c
����*^8"�  @��ƃ"��_,!D�Ǜʌ�9�^����ɏ�����r��-�s��A��cM�����l�J/�I�\Lsa���9$D:&@j"~9�r�O?�YӤ���@)IP&��/a���u���7�.���ŧ�'���4/�J� [��L���8�#��dr�r0 ��T�����b�?�"�m���T'�m���Z���+Tʡ)|熛��2�KNZ���*���r����½;�)��U�\�	��R��w���6�����m�����Vv�&1�0Q ��U��s��	6&����#,)��n�$�oP~�!�O��7��jZW�=�m�NC�R=�|�aD�Ҳ͔V��A����!�z:�yŒ=�*BMq
5%��in(����B���,�A�M=>;W������kZ�������C��8;3�y��ܾ�ˊz�x�>��xO���O�v�UujJ���!&����`!'[,^Ls&hx������S�=M�T��ɿ[����N�����µ�x�RRi�V'I�9+�e�͌=�E��3��F
���Gl1�p' ��8������c�135M�LYO�	�=hƨ�;*q0L�+�[[�=9Us&if�>�H4TXq����F)�sb>*q,mT�8%�M㚀��Z��ċ"r�`�y'�{aX�JoCe컶�-�3�j�
� tt߈��F+��a_B�T}!�����k&gJ���՘7ԥ����Ұ�`}�K_R��!�[e��{���+V�2�5OX�"L��]*�^��XE]~J΍끅�0�gO�J���{kT'��#��^�����C���7@�N�k��Z�cǔq'mz)��FCECU���Y�~���4mj���e�m��}Ki�-a�g ��;Ø�$���y����6��������-�F����Z���wu��I[5��,7
r��o�jV۫4���	���H�5�����Zs��\�7_��,n�E��L��m�aЫ�F@�Q��x��lC����y�٠c=}�Uu%��UE���T�@��U�$�O?��p,����� h��FNB��Ւ)��sF���]yþ�g_�o����羽�TJʟ�u�ۗ����D�Ji��/�~�ŗ�g��O����S/8E���I;���D�H{عO���N~�I���JN�����{9ձy�-�ѩP��0z}c�B�\�'����Y5�S\{Z��w�Ƨ��O,-�M�9�� Jhd(#�D� �D�-䆎I�!����U6�K�ȸu�:oڪ�̣c�ڦT�FO��Ƌ]:@�m �z-�e)����z���CZ��/��ԣf
p�3�c�G�"����f/@�gU��
/�*n�h7�K��JúH��c�Qա�\Sbp VU
CK�V�l2����8��a�� 3�E�sF�� ��S�j��_St��(5���EF�!��Zi�Д���j�s\�ڦ~��견�e�9�"��T�Iu��yƔv^By�$BX��c���kv�p�A��O'3�ㄝե~�y��b�1�_�6T�,7 ��$z��n�i���l�O�~e�U�5�Q�a�ƇB�ŲM����^���	��1/��Q��^,��� o����7|s�QN_O~��F����c�R�Ê&�����ޡ1��{y���utb��S_�޲���ͭ�i
�������U��|����t�0?X$�������+2��j�Wh1�~Ȅ�9���xު��g�d���_qW����v���y��5]���+˦�"쾽����%�"��؍��8EQ������ ����-��z��!�Ŕ�)��@wF�A��94�{KXQ�;�d��|�4���D��X�v�iG뇏 r��Oz2[�:��5.�����c�|o�MD-��-���� �S�@A��I~�u+.@Ct:%%ʞ�f\�WZhKT�b��nl����6�6��BK�r2���8�H8B>˸9rD=�v�:1M�UDGp�b�h��`�UPś{�5,d�����(�g�ki.�P��:T��>[� F*���%P�U�RU����(@���g(�c���|�ۤ�V1���C�C-,X���je��@H{%��q����' կ^Z��ej)�>�ܰY��2���J�6*D�^�T�A���r+�i�<[��T��
f$@m!��ܙ�J�����d�J(iA����տO_G����&��2�(���B5�J5��B��b���T��A��zp���ҿHMdQeD�ٰʘhr���fƟ֕A�+�ܘS�������σE���_Z7��
@�,��3YI )�*�ٹ�ؿ-��F����i�w��G�O�+������+!N�-�A�k���#�-q��r��xV��5<�����X�W�����?�_}��A�AK~]s��o�뾗�T�n*��.�⏓4-�8��R[N6�"Rж�Y2�RKo���=��uq+�T15>\̈$�b��Fqg7��pqX+��	h��%��x�@N;2��]C{X��E�� ����ig`�b�0�\�#7*��J�5?.,̮�Y|��}\/� �[rZ�C>�צ�p�t�^���ߌC*^�
F�B����� X!�kTA�2�H��:pM�ƪ9[m}�R�@�tw2�`pRaJ�pd���Q1t�g�3Tn����tn/iOĖ�M|�Z�H��s<�u�b�J�6��� ��8~��p<g�$p����i��븴1@�C1D�
� )�<o��V�a6�}E��;��V���YZ�G��5.Qp��r�J��r0zV�*+�3)��E�_'���
A���F5���J��lJ����?��Q+e�����r���!��l1^�emK��2��:�J-0��>�k�R6yo�C��R�q��&�gzt����W�a����xhs6!�rZ�gT�V$}��q��B�\.�Jy3����\HC�:�3mVb�.=���� �������E������JuU�3ݧ��$�[(�*��M����+����S��Cݶm��C=��O��t+9�X� uX���Ɇ�ꮆB�Úв�?���$��⟓�������DeY�$�4��b5�bv��-a��3��9�������7���]�e�ڻ�\s�ͯ8�?�����eԤAӀob���!ʴ�܂C?yN;�ű�����Ď?��ݹz���!Z6�}�69�t]���y����
5,_�w�:pց�V�-�
]��\Ӕ �|Hm�v]j��;֟�}���Y�'Υ���]k��|8H�
��~v0�},�g��y��hg���iG@9���M�wB�pjF��ӵ���~;yמ �b����n�B�;��tTa�RlK-�*�8�EH�ȗ�V,@B��¿x�Ƅ�V�/�e�8;'GSQ�����2�o�H:�)\F�M�=��<�7����n-,�{F[�Yo0�:!Qv���>I�!0X�z��dz5��U�M�I�Ka.�Dr�֞B܁k͘��;���a,QdM�AHs|�\3���X,,�Wu�|-�.S;�+f2Y�7����;e�%�MFk�ߌ��|�ar=_��B�+��T�̘=Ӎ�c,��`���){�o���F�0h鹧����ʶ�zN۹������=������{�145�Ue�L�%@�Ҩ�ǌ���������r��zY k��8حu���E3ݣE��M3څV�V��בɀJ��[ղa�����򚳮��ES]�����_���_��\�����K��x��׮PCL�+��gFxh~��>1y�b��>'�P'�5�o���'̲(�~���Y[f����CA'����̼��y^W��b���{4��k�`,�1U�D� �	 �uk��t��g!�>]�O��"0IvJ��9���^i�.FE�LG���X̒�p*骑Up~�0��'�K�!ZoDw�?�N��M/�e�gEd ��S[l�yh׶p��lҌY�Z��b�B�@��V#��j�n[;増�� :���.lLX}'}���(7�V�3���^�Z3{1�gi���EGz�v�@� ô�ƗIS5)V�O�g���x!'��<��&�h�QUSzLN�z�Emw��	�`��h�Q��a�k�u�����J����y�9�����|�,}:eFZF �$��6�`1���,;^6>���2��g(6�5���1d-<sșw\[�>��X՟��q��8�L��æ�ã�&�/.)k��~��;���3�n�rP~�ׁљ��~��'޳�೫�V��S�ƼBe�T@�ácG�7/�o�M�3\z����2Z������X��G���ytY��9��,�J�],]�K�J�^|���g�5U���������M��SG�u�����54�M55��ssǏw�t�l���笽{�?������w�l@vgM���H���h/,;)��Ӓ{�4go��W�����ŋvJ�~(L�bg��XŬ���s<�hXp�񓛵�t��Y��9�3ӑD���ȼ������o�-Td�X����T,E�8N��� �A�t�'j~ _�1�/c�����7{*�Y��Tw�.���5���޿�� Qr�&D��*�}�0^z�J��UV���5c�5�k�� �]+���X'�������?k M�VvarıכP��Ҳ����R�{
eΉ���9����P ���P��k?Q~�F���ʂ�E��ήcV!��vu�`y�4:z��A/Ay0N{�c���I{����%���Wl� �;$�n�FJ��r�%���TBB�SXbY�X��DB:�$����}~ߞO�aΙ3sf�+E�D.����^U���b�h0j�E�K}�H�dW~��Dz)� V��&�W�i�%W���D	X�����8�j'����n5Or���W��em=�l��#HD�����`��Z§�)cs����L4Ϳ�>�33zݝ�F�z�?z��^q��'��YX9��~�<�+���g��+����g-�7�?n5�յj���ZV�z���&4n	(e�.�/f46�P���;������:Z+�`�O��}���5j�a��͍���8��c�,)����=����yj��2Z�6�٫��	�S,�I��N#�`���?�Cc�k޷���c
��%5�?�)#Qy6�y%��1��ʼ��+�]�|hE���s��07r̀�v:��v�Z��Y�~M�{c�X����Q%�}��T��o�$rrs�L#"�<B�49Y[Sa�[a�J{�̾��tܖ?j�B�����v��w�4WLb���-B�ؠ��Z���8[B��7�+�W)y�O♇vE�?=x��u�SQ���wLS�����ڥ|��kK��C25���1��V�x�}$�>>��&�Y��� ���>%�t�䩪�����Bz���W?/�.U7c5�y�ꁶ����^*�Ӱ ��'�R��8%�ت`D�A4�c���jQ W)�l6V���O�=|J3mbH��J������n��}U<>����y�W��)����6�2ʃ'���K�d�'��y��y�iH��-�J�e�^K���DK���[��v����m�mAJ�jb�\����Wb�_*z�8/�/:#�C��J�>f����e��"Ҿ��4LKy��?��i���I���l�9!�q��u/�g�}����x�7�I&����w�KKjƟɴ�A��_�Ǒd?-B��BT�W�0�b�s���\=S���2dh��"�?c�ޓ���w�Ŋ�u�7k��1>�+�=�0�w�x)�g~`��Ӊ^3h@ ��#�­C(ͭN����E����p@�V�҂/�����d%�|x���Qՠ;�M��V���ff���1Nǆϐ	��L��mEѮ�}�#����s2�񿞲���X8����h�"*l��UcݽN�T~���ZwدS�柤H+���4<�4ܶ%xG�V�ݙ�9k���>�0ҙ�\���B�pS8?��3Vh��*�G&,iL���C��!��Ɉªҙ�|H���K���t�74���*�b�{2��$�&��e����[ǳ�1G�8ô9�� ϔ0F���]9��q"l��ʍ�mZ��ԥ�ta��C��3��1r����*T�Ÿ�T��3��ۮW�q�Ue��J*@�L��u@a���?�?�/�rj���y����i{>�/ڮ���q~_۠�'b칀|�-��:��v��-&��ۂ�-�'��R�4U�u�U�Y�݈�SАbI2m.��)~B3~��̰v��f~���0}��in3l��C8^�Ig����j ��
���`���7x�d��&NHdR9p��C}J'<U��4�_�O�ŴO�)����"���y�4j�P���3B="�;^�����Z}��-�г���t9�j*�@6P5$�lkrx ��e0ԡe�v0���.ݶ.��8}�&�>�k(�~u�03�=��h����e>w�����_�������L�>�8�q������k�F�G�]je/w�u���W��:����]�S�>�:�;��՝L�^\�m��'�"��E��c��Ɋ�D����UH�h���k��FGKw����$8w0޷� K��n�f���wR�*����!���M�\��o��Y�+y�=C���}����l<g�F�p2"�k )s(���ɠ'��?G����I6��O�7��*֠�3�bo����rJm����@kr ��M�-���9����jW�`��āT����.�d��UD ���Ф*�_�uW���9�3����ΒP����4�%���/7Љ���Zܤ.��C�Wk�[����TC|˥���:�6�њc�͍]����u#\c�$,��ت_�ϸ��r�����;���*������ ���cs�U�[Y1%oO1�4�� U�5n�6΄A ���Q�^�f����;U4)�y݁�\@#c�B�8�z$�H���:F6BX����#3]�/�m�A����Z{�M~j¥�|g7�߼�qqfC`[N6��}]�f_��}�$��g�\Q��n�T�d	9����&�����6z�b�V�_l���fJ���E	��ӑ9d����l���M�s�;�|���9���MY;4�-]Uo|��t���@���<��ĭr�op-�_4���1����-�ű1P
�5 ��(�\�j�W�n�>��������ۅ�eJ���2�����[cg�_��
�L^n?<�xY���� ���{�ۍb�k .�>MZ�����\:]��z:�X�%�B~fwX�
:\6���M~���m��H�������suC2j!�����`������vf�6��+��b�ū�=%J�ˑ�2DDR�����|5�㸐^Y|x��VܟL���~�&/�ˋi�����@� گ�{����K�
Vh��bDG��Ƥ�<�H��%G<*:i�Ax�0L�K��̊��_����x59�������N�?1�Z��1�$��M���{�P�x���E����RGJ��;����*{�M��lh,�ᙅA����`��)����c���1lD9q�'�+1F)�Lou$|Ø�	(s�N.�_���,�v������oh�MPT_�W
C� �oUǭ�k�Jڤ翵�ɾ�ƫ!���F��G���Dsهsc��J��Ĭ�F�!֫�L��?��Xvw�z��d�$2J�s�#4�Mc�˸g���H1�����=U��|���Ϩ�g��g��]f��=����5�!�f�FD��"M��&��_�������)�E��%��G�RO^���7p}ǽ���*���w�A���\ķr��G�Z�u�<kz3@�TjS�<�K��}�Zj��v��^�2H�Y�"٪hg��n�|�&I��^�OF������$dd���,S(q�W�f0�f����Ӗ���U����9�6Iw4vW>`�c*J�f_�g��{&��t_���]z��q���|����/��Fv�٘�r�v��9�ڄ��S8��-����y�*VV�+��f�6ᕮ��M�l��	JB�t,|Et,��Lu���$�&�}-�r��M��6 P=�G�ԏ��X]��^U��	��c�+�C!P�r��Zs�ċ!��̫ -�9�}��-�m�[�PT:cM�z��UnV%��Vs�j\$06��V�M��}��Ķ%��!�5������<
��K	�c7t������������̤�ͫ(����''�T� _P����\Ca��Y�,N�*jU�L4{��Du�Yw�'����|y�o;�`�?�,,��_ʌ�RHWb�',���֢g��=����2������34���p��'�s����F��²�'>y�ա��f�7���,.��B�����0�]�zM@��It�w�iM�u�l2ι۹����WM{H�S��Ÿɹ"��[0-׊7;}�9*|q
��y����	�|����ͤ,41��P~��z���il_�њ?u�Q���ף�9��5׼' �%p1�\��`t�����%�W���D����H���Vs#���2����dJ]���޸j{6�Y֟�ӱ�38�N�J�,�$���٩5���q5�������5 9d�I�Z~A}�m�<7v^=&���F�f-���(kMuS�O��>�yW�Eb�i��ix��W��kL�*�$`�x�ko����V��㴑����l�J�"
�X�����9B�����{o��;���b�m0��s16���+5[K��r��]�0�Y�/h,����I�q�H��-[5l_iQ;C5�����2��o/�_	`>�'o;e���|k KX����[KiB%�/���V^qX>O@.W���A~"�x� �k�4"]����N�$\������Y���<;f���^)�vh?�OΙ�0�((�O����&���*�H�=��Nw�}F�_��%���İJ�,��шw۬|3���g.�/g`9(��&&���sB��OK�q��G�k�U$A�-����ь��X�Ix�V=�cNq!���� /���gt���E0���]Ll�k���AO �R&'MyvG�Y��������ӅnR:97�o:�\�+7J�d����.���������%ϩ���sf�ԗ/��Ņ]����>I%N5z;�p��g�^#�"����dl4�C�2���[]6?Ȑ�/M"��;���!����ǉ�']hK-&@��d�V�Zt��x_K\��lΊ�%��'��m���o���8�K%��<���]���O΃��O�ϯa:�Dr����О�� ��3.�u��R��}j���	t
��^�gSD���||����c�Pi ��-E������MDF������)#Щ��'��e�ֻ3E�K�o{~� 敜TU��]�?����&<��1��g����NW%<g5��.4J��rx eX��pB̮�cl,{2j�}�6��q�b�'��n�a��� �Hc��� ��"y��>I�(�=4,i����>�>��;�&^��B�I�]����IKt �:B-�b�Q�F�@�\�Nm^�3�2�v�\��ⲵ�r�bY��L���"Ĉbc��1���a�0�J�iP��[��Y52q��
"	~��F�1fNk��v~lI�)Vc���^�~G�����3�*ԝ���&B��3���O��}��-�����"W���Ե��Sxc�d�X��X?J�my[������L���@,�_�V����QZ�Ca�n<�EM�A���1�p�k�f��� {�h*/uٲ-���v�����Y�㷫�	���ʟ������J)�s(�v1��1�8��}G�7�cs<ǎW���u4����9CC��ᓷFji��$�i	D^T�o�mx�}��٦7�-���99#�ΤN��z5�Y�D����4�E~�F�獓S������۩�#F
��.��;v�:ԓW=H7��Yç�Z���|�l���4�l�a;2���m3��tcɗ 5��I��HHE(S���eγY���Z����ji��RV�m�ZezY\��k$� �];�#z-����!!%���_���<��g4=U���<���E����;�D+F-~[��t4��u�b�0\��amַ̀���tS�2TJ�U�uehٵ�(�Kj�J'g�vlQ�}]��U�#��x��N��d,��G>�y̡(��㰞p ��4���!�2��AA������(kp2��	���ک�е�
�X��F�6Ū�_"M�
�91!�h�)�Q�hb��ph��6 !!~�Go�i��p�/�@����>�A�n�=�u:�8��pK�0W�4�n�K����q`e	wW�;��?ET�c���q���6��a,d�.CZq�/tX� ��ϼ�%J������O�Kͷ��/�Wx] j��,�MUjB���ZtV� �SLo o��11�P����fO�D6���h�i�3�b��I'	f'f���ct���������R�������N��6/O\\<nI<q����&�Xh%G�グ��z7ҁYyS<���hbcE�jû�[)i�ގ�+tusc��4	

j�+�GP��@x��a��|��eֆ)Х[oS�k~��;0j?�T�c��iy�u����xe;{��j?Z���B�-='�ɟ�!󷓯�\��ke�
er�������:յ�ňm���p� �0���i�#ڱ6��6qO�����(�X�5���C{	�n��)V���A+�Wɛ6��!D�)�u)��Y�E��/�	҉)�������a2������V�Id���5zvV:�c�.��ݵ���@��27����XK�&$m���_��/�Z�����?����[����,sN�ti�J%�OSUO�^���� PK   �
.X5	�cm  �%     jsons/user_defined.json��ko�6���`죩�~ɷ�Άl�v��A��V�+y�$H���QIcy���P����P���C��`������nc�vQV�wv�)��]�)N��e��7�n'}��e��y��"!��%<�����ݟg[��^?��3<��i8(�T��Vs͐�"�	As�
d
)*cs�	��ˣ'����2��|]����l�x]������[��y��'����ܬ��è^�wP�RI8s���&�}s�����s���U�?;7�꼘nץ�聆��ޔ�H/�e��*ťlT*�R�]��ʿ�k����.��m����q��>�	�_d��`|~�>�nG� �����x���i1n�U}_��l�O�ze���I����I3���^�&��G��Ѥ�UE2�����z��dl�2̑P#.�2����Y̕"v>?B������
L�O��b�/$K%7O��8e3�/7��'|������z	���q���i2����Ur]�;�Lw���!�����B$�H�l�ad��3_�7�(�sep΄������HJ�X*���j�EJ��n8NY*� �_Q�1y��W��6FZ-H� ȗ���� �Co�
@�mLf�-�	ϩ�	s�+�K�`R z
xW� k�k�YU6��l�KY%�e����J+�Xd	S�B�6R!e)�'=m�f����˔(n�fvרT�ě�a�
�RΈ[U�i������A|��J5����(�З%�&> �+�.o�&�m!� !��Md׾�54�(޼`�w�{]�ou�q����2,�\,�V8T��hn��Z�=O��VS�!�!%�M;5�{�9�]��I�B�)W�~��I�s�!�%�Q���#G�\��ܕ��ؕU��ܟ	���F\9��?�R��)#3m&jqԞ��Yʔ���k�i^��&.��8Uj�o��ɟ1i^���R�M���BD�4&�s`1��x�O1)��x�����x�T7��J_T�� �[�t`|��x�	�s��,�������;$�����+`ш�����߱$�hҵ��Vm�  Do!h�[!N'g?�]_��u�B���i�u6\�C�~#��>HM�4Q=��z�QcbaSPO�v��X@��S����A=UZ��5���D=���ˀ!�C�����f?U.UA ���������ھ	,}�_���v�M�hU�A�����&���mf�~�`�f�&��m�.��%�����m��OZ�4��D��m�x�:�<e�`��[�[���~�nϚV毧��5�5x�؄ ~}����(��=�u���%�E���ZB�Jy��E^8�`H�y��p�ceAz�	pe,5�h�;�\�<�
&R���J�T�x����C���t�꭭ܨ�Z����r�ɭ@�q���X �#+e�c�
���5թ�\{{Ǆ��i,�/���>!���/6���(���[�_倫�����nu����=.�
z>V�%W�MF_2g�e2�n�`�QMq��4���"�L���6�R���= �!�Q�rl�7��T�=�&�I��r����Thb�h��t�=%v��@�Η������-��^�ӧ���&/�0~��Ͼ��ρ��҂�@�0 ��
�w�����/PK
   �
.Xƨ�mL  1�                   cirkitFile.jsonPK
   �-X����%a 3c /             y  images/26e5b11e-e137-4512-8967-7e228f6738e0.pngPK
   �cW�����8 �I /             �x images/31d687a0-e383-4fc9-9100-a6b790c355a8.pngPK
   WL� �� �� /             � images/3344f319-942e-4277-a6d0-796a8e5017f8.pngPK
   M��W�&
�G_ �h /             ��
 images/56c78dca-afcd-4253-86bc-452069e6d2d2.pngPK
   Ԣ�W�@͎� �� /             N� images/633b3a04-5760-46d4-a0cc-eb31fb771ebb.pngPK
   �	.X�:sJ� j /             )� images/920576d2-9ce5-4348-9cff-973310077ed8.pngPK
   �-XS��
�M 2T /             � images/a053b5f3-ee57-4c4b-b9e3-486563af4e78.pngPK
   :�-X�L�,� o� /             �F images/a0820d33-a834-4c8e-839c-8eeec59e25c5.pngPK
   �cW���/�� Z� /             l images/d3087b83-655e-4811-b17d-9d66f7a3b2a5.pngPK
   �
.X5	�cm  �%               Z� jsons/user_defined.jsonPK      �  ��   